magic
tech scmos
timestamp 1700198425
<< nwell >>
rect -326 1 -224 22
rect -149 2 -47 23
rect -301 -90 -265 -71
rect -258 -90 -231 -71
rect -115 -84 -79 -65
rect -72 -84 -45 -65
rect 16 -77 63 -58
rect 72 -77 99 -58
<< ntransistor >>
rect -315 -23 -313 -18
rect -289 -23 -287 -18
rect -264 -23 -262 -18
rect -238 -23 -236 -18
rect -138 -22 -136 -17
rect -112 -22 -110 -17
rect -87 -22 -85 -17
rect -61 -22 -59 -17
rect -103 -108 -101 -103
rect -94 -108 -92 -103
rect -289 -114 -287 -109
rect -280 -114 -278 -109
rect -247 -114 -245 -109
rect -61 -108 -59 -103
rect 27 -109 29 -104
rect 37 -109 39 -104
rect 83 -109 85 -104
<< ptransistor >>
rect -315 8 -313 13
rect -289 8 -287 13
rect -264 8 -262 13
rect -238 8 -236 13
rect -138 9 -136 14
rect -112 9 -110 14
rect -87 9 -85 14
rect -61 9 -59 14
rect -289 -83 -287 -78
rect -280 -83 -278 -78
rect -247 -83 -245 -78
rect -103 -77 -101 -72
rect -94 -77 -92 -72
rect 27 -70 29 -65
rect 37 -70 39 -65
rect -61 -77 -59 -72
rect 83 -70 85 -65
<< ndiffusion >>
rect -316 -22 -315 -18
rect -320 -23 -315 -22
rect -313 -22 -311 -18
rect -313 -23 -307 -22
rect -290 -22 -289 -18
rect -294 -23 -289 -22
rect -287 -22 -285 -18
rect -287 -23 -281 -22
rect -269 -19 -264 -18
rect -265 -23 -264 -19
rect -262 -22 -259 -18
rect -262 -23 -255 -22
rect -244 -19 -238 -18
rect -240 -23 -238 -19
rect -236 -22 -235 -18
rect -236 -23 -231 -22
rect -139 -21 -138 -17
rect -143 -22 -138 -21
rect -136 -21 -134 -17
rect -136 -22 -130 -21
rect -113 -21 -112 -17
rect -117 -22 -112 -21
rect -110 -21 -108 -17
rect -110 -22 -104 -21
rect -92 -18 -87 -17
rect -88 -22 -87 -18
rect -85 -21 -82 -17
rect -85 -22 -78 -21
rect -67 -18 -61 -17
rect -63 -22 -61 -18
rect -59 -21 -58 -17
rect -59 -22 -54 -21
rect -108 -104 -103 -103
rect -104 -108 -103 -104
rect -101 -108 -94 -103
rect -92 -107 -90 -103
rect -92 -108 -86 -107
rect -66 -105 -61 -103
rect -294 -110 -289 -109
rect -290 -114 -289 -110
rect -287 -114 -280 -109
rect -278 -113 -276 -109
rect -278 -114 -272 -113
rect -252 -111 -247 -109
rect -248 -114 -247 -111
rect -245 -112 -242 -109
rect -62 -108 -61 -105
rect -59 -106 -56 -103
rect -59 -108 -52 -106
rect -245 -114 -238 -112
rect 22 -105 27 -104
rect 26 -109 27 -105
rect 29 -107 32 -104
rect 36 -107 37 -104
rect 29 -109 37 -107
rect 39 -108 45 -104
rect 49 -108 57 -104
rect 39 -109 57 -108
rect 78 -106 83 -104
rect 82 -109 83 -106
rect 85 -107 88 -104
rect 85 -109 92 -107
<< pdiffusion >>
rect -320 12 -315 13
rect -316 8 -315 12
rect -313 12 -307 13
rect -313 8 -311 12
rect -294 12 -289 13
rect -290 8 -289 12
rect -287 12 -281 13
rect -287 8 -285 12
rect -265 9 -264 13
rect -269 8 -264 9
rect -262 12 -255 13
rect -262 8 -259 12
rect -240 10 -238 13
rect -244 8 -238 10
rect -236 12 -231 13
rect -236 8 -235 12
rect -143 13 -138 14
rect -139 9 -138 13
rect -136 13 -130 14
rect -136 9 -134 13
rect -117 13 -112 14
rect -113 9 -112 13
rect -110 13 -104 14
rect -110 9 -108 13
rect -88 10 -87 14
rect -92 9 -87 10
rect -85 13 -78 14
rect -85 9 -82 13
rect -63 11 -61 14
rect -67 9 -61 11
rect -59 13 -54 14
rect -59 9 -58 13
rect -290 -81 -289 -78
rect -294 -83 -289 -81
rect -287 -80 -280 -78
rect -287 -83 -285 -80
rect -281 -83 -280 -80
rect -278 -81 -276 -78
rect -278 -83 -272 -81
rect -248 -81 -247 -78
rect -252 -83 -247 -81
rect -245 -82 -242 -78
rect -245 -83 -238 -82
rect 26 -68 27 -65
rect -104 -75 -103 -72
rect -108 -77 -103 -75
rect -101 -74 -94 -72
rect -101 -77 -99 -74
rect -95 -77 -94 -74
rect -92 -75 -90 -72
rect -92 -77 -86 -75
rect 22 -70 27 -68
rect 29 -70 37 -65
rect 39 -67 57 -65
rect 39 -70 45 -67
rect -62 -75 -61 -72
rect -66 -77 -61 -75
rect -59 -76 -56 -72
rect -59 -77 -52 -76
rect 49 -70 57 -67
rect 82 -68 83 -65
rect 78 -70 83 -68
rect 85 -69 88 -65
rect 85 -70 92 -69
<< ndcontact >>
rect -320 -22 -316 -18
rect -311 -22 -307 -18
rect -294 -22 -290 -18
rect -285 -22 -281 -18
rect -269 -23 -265 -19
rect -259 -22 -255 -18
rect -244 -23 -240 -19
rect -235 -22 -231 -18
rect -143 -21 -139 -17
rect -134 -21 -130 -17
rect -117 -21 -113 -17
rect -108 -21 -104 -17
rect -92 -22 -88 -18
rect -82 -21 -78 -17
rect -67 -22 -63 -18
rect -58 -21 -54 -17
rect -108 -108 -104 -104
rect -90 -107 -86 -103
rect -294 -114 -290 -110
rect -276 -113 -272 -109
rect -252 -115 -248 -111
rect -242 -112 -238 -108
rect -66 -109 -62 -105
rect -56 -106 -52 -102
rect 22 -109 26 -105
rect 32 -107 36 -103
rect 45 -108 49 -104
rect 78 -110 82 -106
rect 88 -107 92 -103
<< pdcontact >>
rect -320 8 -316 12
rect -311 8 -307 12
rect -294 8 -290 12
rect -285 8 -281 12
rect -269 9 -265 13
rect -259 8 -255 12
rect -244 10 -240 14
rect -235 8 -231 12
rect -143 9 -139 13
rect -134 9 -130 13
rect -117 9 -113 13
rect -108 9 -104 13
rect -92 10 -88 14
rect -82 9 -78 13
rect -67 11 -63 15
rect -58 9 -54 13
rect -294 -81 -290 -77
rect -285 -84 -281 -80
rect -276 -81 -272 -77
rect -252 -81 -248 -77
rect -242 -82 -238 -78
rect 22 -68 26 -64
rect -108 -75 -104 -71
rect -99 -78 -95 -74
rect -90 -75 -86 -71
rect -66 -75 -62 -71
rect -56 -76 -52 -72
rect 45 -71 49 -67
rect 78 -68 82 -64
rect 88 -69 92 -65
<< polysilicon >>
rect -73 50 -27 53
rect -295 44 -193 47
rect -295 34 -292 44
rect -264 34 -206 37
rect -330 23 -287 25
rect -330 -33 -328 23
rect -315 13 -313 18
rect -289 13 -287 23
rect -264 13 -262 34
rect -238 13 -236 17
rect -315 -1 -313 8
rect -289 5 -287 8
rect -315 -3 -287 -1
rect -315 -18 -313 -15
rect -289 -18 -287 -3
rect -264 -4 -262 8
rect -264 -18 -262 -8
rect -238 -18 -236 8
rect -228 -6 -222 -4
rect -315 -33 -313 -23
rect -330 -35 -313 -33
rect -315 -40 -313 -35
rect -289 -34 -287 -23
rect -264 -26 -262 -23
rect -289 -36 -283 -34
rect -238 -34 -236 -23
rect -279 -36 -236 -34
rect -224 -40 -222 -6
rect -315 -42 -222 -40
rect -209 -65 -206 34
rect -122 34 -119 49
rect -153 24 -110 26
rect -153 -32 -151 24
rect -138 14 -136 19
rect -112 14 -110 24
rect -87 14 -85 17
rect -138 0 -136 9
rect -112 6 -110 9
rect -87 0 -85 9
rect -73 0 -70 50
rect -61 14 -59 18
rect -138 -2 -110 0
rect -138 -17 -136 -14
rect -112 -17 -110 -2
rect -87 -2 -70 0
rect -87 -3 -85 -2
rect -87 -17 -85 -7
rect -61 -17 -59 9
rect -51 -5 -45 -3
rect -138 -32 -136 -22
rect -153 -34 -136 -32
rect -138 -39 -136 -34
rect -112 -33 -110 -22
rect -87 -25 -85 -22
rect -112 -35 -90 -33
rect -61 -33 -59 -22
rect -86 -35 -59 -33
rect -47 -39 -45 -5
rect -138 -41 -45 -39
rect -31 -51 -27 50
rect -320 -68 -206 -65
rect -131 -54 -27 -51
rect -320 -94 -317 -68
rect -289 -78 -287 -75
rect -280 -78 -278 -75
rect -289 -94 -287 -83
rect -247 -78 -245 -75
rect -320 -97 -287 -94
rect -289 -109 -287 -97
rect -280 -102 -278 -83
rect -247 -94 -245 -83
rect -131 -88 -128 -54
rect 27 -65 29 -62
rect 37 -65 39 -62
rect -103 -72 -101 -69
rect -94 -72 -92 -69
rect -103 -88 -101 -77
rect -61 -72 -59 -69
rect -131 -91 -101 -88
rect -246 -98 -245 -94
rect -279 -106 -278 -102
rect -280 -109 -278 -106
rect -247 -109 -245 -98
rect -103 -103 -101 -91
rect -94 -96 -92 -77
rect -61 -88 -59 -77
rect -93 -100 -92 -96
rect -94 -103 -92 -100
rect -61 -103 -59 -92
rect -289 -117 -287 -114
rect -280 -117 -278 -114
rect -103 -111 -101 -108
rect -94 -111 -92 -108
rect -61 -111 -59 -108
rect -247 -117 -245 -114
rect 7 -131 11 -85
rect 27 -90 29 -70
rect 37 -81 39 -70
rect 83 -65 85 -62
rect 27 -104 29 -94
rect 37 -104 39 -85
rect 83 -89 85 -70
rect 84 -93 85 -89
rect 83 -104 85 -93
rect 27 -112 29 -109
rect 37 -112 39 -109
rect 83 -112 85 -109
rect -207 -135 11 -131
<< polycontact >>
rect -193 44 -189 48
rect -296 29 -292 34
rect -266 -8 -262 -4
rect -232 -7 -228 -3
rect -283 -36 -279 -32
rect -122 30 -118 34
rect -89 -7 -85 -3
rect -55 -6 -51 -2
rect -90 -35 -86 -31
rect -250 -98 -246 -94
rect -283 -106 -279 -102
rect -64 -92 -59 -88
rect -97 -100 -93 -96
rect 7 -85 12 -81
rect -214 -136 -207 -130
rect 34 -85 39 -81
rect 24 -94 29 -90
rect 80 -93 84 -89
<< metal1 >>
rect -320 37 -273 41
rect -320 12 -316 37
rect -320 -18 -316 8
rect -311 29 -296 33
rect -292 29 -281 33
rect -311 12 -307 29
rect -285 12 -281 29
rect -311 -18 -307 8
rect -294 -18 -290 8
rect -285 -18 -281 8
rect -277 -4 -273 37
rect -269 24 -252 28
rect -246 24 -240 28
rect -269 13 -265 24
rect -244 14 -240 24
rect -277 -8 -266 -4
rect -259 -12 -255 8
rect -277 -16 -255 -12
rect -294 -25 -290 -22
rect -277 -25 -273 -16
rect -259 -18 -255 -16
rect -294 -29 -273 -25
rect -235 -3 -231 8
rect -235 -7 -232 -3
rect -235 -18 -231 -7
rect -269 -27 -266 -23
rect -269 -30 -251 -27
rect -243 -27 -240 -23
rect -246 -30 -240 -27
rect -283 -56 -280 -36
rect -193 -46 -189 44
rect -143 38 -96 42
rect -143 13 -139 38
rect -143 -17 -139 9
rect -134 30 -122 34
rect -118 30 -104 34
rect -134 13 -130 30
rect -108 13 -104 30
rect -134 -17 -130 9
rect -117 -17 -113 9
rect -108 -17 -104 9
rect -100 -3 -96 38
rect -92 25 -86 29
rect -80 25 -63 29
rect -92 14 -88 25
rect -67 15 -63 25
rect -100 -7 -89 -3
rect -82 -11 -78 9
rect -100 -15 -78 -11
rect -117 -24 -113 -21
rect -100 -24 -96 -15
rect -82 -17 -78 -15
rect -117 -28 -96 -24
rect -58 -2 -54 9
rect -58 -6 -55 -2
rect -58 -17 -54 -6
rect -92 -25 -88 -22
rect -92 -28 -80 -25
rect -67 -25 -63 -22
rect -75 -28 -63 -25
rect -90 -46 -87 -35
rect -193 -49 -87 -46
rect -334 -60 -280 -56
rect -334 -103 -331 -60
rect -301 -74 -264 -71
rect -259 -74 -231 -71
rect -294 -77 -290 -74
rect -276 -77 -272 -74
rect -252 -77 -248 -74
rect -285 -94 -281 -84
rect -242 -94 -238 -82
rect -285 -98 -250 -94
rect -242 -95 -229 -94
rect -242 -98 -210 -95
rect -295 -103 -283 -102
rect -334 -106 -283 -103
rect -276 -109 -272 -98
rect -242 -108 -238 -98
rect -233 -99 -210 -98
rect -294 -118 -290 -114
rect -252 -118 -248 -115
rect -298 -121 -239 -118
rect -213 -130 -210 -99
rect -174 -97 -171 -49
rect 17 -61 63 -58
rect 69 -61 96 -58
rect -110 -68 -72 -65
rect 22 -64 26 -61
rect -67 -68 -45 -65
rect 78 -64 82 -61
rect -108 -71 -104 -68
rect -90 -71 -86 -68
rect -66 -71 -62 -68
rect -99 -88 -95 -78
rect -56 -88 -52 -76
rect 12 -85 34 -82
rect -99 -92 -64 -88
rect -56 -89 -7 -88
rect 45 -89 49 -71
rect 88 -89 92 -69
rect -56 -90 4 -89
rect -56 -92 24 -90
rect -111 -97 -97 -96
rect -174 -100 -97 -97
rect -90 -103 -86 -92
rect -56 -102 -52 -92
rect -10 -93 24 -92
rect 2 -94 24 -93
rect 32 -93 80 -89
rect 88 -93 96 -89
rect -108 -112 -104 -108
rect 32 -103 36 -93
rect -112 -115 -74 -112
rect -66 -112 -62 -109
rect 88 -103 92 -93
rect -69 -115 -51 -112
rect 22 -113 26 -109
rect 45 -113 49 -108
rect 17 -116 60 -113
rect 78 -113 82 -110
rect 66 -116 96 -113
<< m2contact >>
rect -252 24 -246 30
rect -251 -31 -246 -26
rect -86 25 -80 31
rect -80 -29 -75 -24
rect -264 -74 -259 -69
rect -239 -122 -233 -117
rect 63 -61 69 -55
rect -115 -68 -110 -63
rect -72 -68 -67 -63
rect -74 -117 -69 -111
rect 60 -117 66 -112
<< metal2 >>
rect -346 69 91 74
rect -345 50 -340 69
rect -345 -50 -342 50
rect -251 30 -247 69
rect -85 31 -81 69
rect -12 46 -5 69
rect -345 -53 -259 -50
rect -264 -69 -259 -53
rect -250 -53 -246 -31
rect -80 -42 -77 -29
rect -154 -45 -77 -42
rect -250 -57 -198 -53
rect -244 -121 -239 -118
rect -239 -164 -235 -122
rect -201 -164 -198 -57
rect -154 -164 -150 -45
rect -11 -55 -5 46
rect -115 -58 -5 -55
rect 63 -55 68 69
rect -115 -59 -77 -58
rect -115 -63 -112 -59
rect -72 -63 -68 -58
rect -72 -124 -69 -117
rect -72 -128 -48 -124
rect -53 -164 -48 -128
rect 60 -164 64 -117
rect -341 -169 93 -164
rect -201 -170 -198 -169
<< end >>
