magic
tech scmos
timestamp 1700324991
<< nwell >>
rect 401 -51 518 -28
rect 159 -105 184 -86
rect 851 -101 940 -80
rect 532 -151 635 -128
rect 161 -171 186 -152
rect 670 -189 761 -166
rect 164 -238 189 -219
rect 799 -230 872 -209
rect 164 -305 189 -286
rect 182 -410 207 -391
rect 81 -450 172 -427
rect 184 -571 209 -552
rect 83 -611 174 -588
rect 779 -625 882 -602
rect 183 -725 208 -706
rect 82 -765 173 -742
rect 183 -873 208 -854
rect 842 -881 931 -860
rect 82 -913 173 -890
rect 616 -940 733 -917
rect 159 -1000 184 -981
rect 484 -1024 587 -1001
rect 161 -1066 186 -1047
rect 343 -1099 434 -1076
rect 164 -1133 189 -1114
rect 248 -1174 321 -1153
rect 164 -1200 189 -1181
<< ntransistor >>
rect 416 -80 418 -70
rect 431 -80 433 -70
rect 446 -80 448 -70
rect 461 -80 463 -70
rect 475 -80 477 -70
rect 501 -80 503 -70
rect 170 -123 172 -119
rect 865 -125 867 -118
rect 877 -125 879 -118
rect 892 -125 894 -118
rect 902 -125 904 -118
rect 925 -125 927 -118
rect 547 -180 549 -170
rect 562 -180 564 -170
rect 582 -180 584 -170
rect 592 -180 594 -170
rect 618 -180 620 -170
rect 172 -189 174 -185
rect 175 -256 177 -252
rect 175 -323 177 -319
rect 193 -428 195 -424
rect 93 -472 95 -467
rect 112 -472 114 -467
rect 137 -472 139 -467
rect 156 -472 158 -467
rect 195 -589 197 -585
rect 95 -633 97 -628
rect 114 -633 116 -628
rect 139 -633 141 -628
rect 158 -633 160 -628
rect 685 -218 687 -208
rect 700 -218 702 -208
rect 720 -218 722 -208
rect 744 -218 746 -208
rect 858 -246 860 -242
rect 811 -253 813 -246
rect 832 -253 834 -246
rect 794 -654 796 -644
rect 809 -654 811 -644
rect 829 -654 831 -644
rect 839 -654 841 -644
rect 865 -654 867 -644
rect 194 -743 196 -739
rect 94 -787 96 -782
rect 113 -787 115 -782
rect 138 -787 140 -782
rect 157 -787 159 -782
rect 194 -891 196 -887
rect 856 -905 858 -898
rect 868 -905 870 -898
rect 883 -905 885 -898
rect 893 -905 895 -898
rect 916 -905 918 -898
rect 94 -935 96 -930
rect 113 -935 115 -930
rect 138 -935 140 -930
rect 157 -935 159 -930
rect 631 -969 633 -959
rect 646 -969 648 -959
rect 661 -969 663 -959
rect 676 -969 678 -959
rect 690 -969 692 -959
rect 716 -969 718 -959
rect 170 -1018 172 -1014
rect 499 -1053 501 -1043
rect 514 -1053 516 -1043
rect 534 -1053 536 -1043
rect 544 -1053 546 -1043
rect 570 -1053 572 -1043
rect 172 -1084 174 -1080
rect 358 -1128 360 -1118
rect 373 -1128 375 -1118
rect 393 -1128 395 -1118
rect 417 -1128 419 -1118
rect 175 -1151 177 -1147
rect 307 -1190 309 -1186
rect 260 -1197 262 -1190
rect 281 -1197 283 -1190
rect 175 -1218 177 -1214
<< ptransistor >>
rect 416 -45 418 -35
rect 431 -45 433 -35
rect 446 -45 448 -35
rect 461 -45 463 -35
rect 475 -45 477 -35
rect 501 -45 503 -35
rect 170 -99 172 -95
rect 547 -145 549 -135
rect 562 -145 564 -135
rect 582 -145 584 -135
rect 592 -145 594 -135
rect 618 -145 620 -135
rect 865 -95 867 -88
rect 877 -95 879 -88
rect 892 -95 894 -88
rect 902 -95 904 -88
rect 925 -95 927 -88
rect 172 -165 174 -161
rect 175 -232 177 -228
rect 175 -299 177 -295
rect 193 -404 195 -400
rect 93 -441 95 -436
rect 112 -441 114 -436
rect 137 -441 139 -436
rect 156 -441 158 -436
rect 195 -565 197 -561
rect 95 -602 97 -597
rect 114 -602 116 -597
rect 139 -602 141 -597
rect 158 -602 160 -597
rect 685 -183 687 -173
rect 700 -183 702 -173
rect 720 -183 722 -173
rect 744 -183 746 -173
rect 811 -223 813 -218
rect 832 -223 834 -218
rect 858 -222 860 -218
rect 794 -619 796 -609
rect 809 -619 811 -609
rect 829 -619 831 -609
rect 839 -619 841 -609
rect 865 -619 867 -609
rect 194 -719 196 -715
rect 94 -756 96 -751
rect 113 -756 115 -751
rect 138 -756 140 -751
rect 157 -756 159 -751
rect 194 -867 196 -863
rect 856 -875 858 -868
rect 868 -875 870 -868
rect 883 -875 885 -868
rect 893 -875 895 -868
rect 916 -875 918 -868
rect 94 -904 96 -899
rect 113 -904 115 -899
rect 138 -904 140 -899
rect 157 -904 159 -899
rect 631 -934 633 -924
rect 646 -934 648 -924
rect 661 -934 663 -924
rect 676 -934 678 -924
rect 690 -934 692 -924
rect 716 -934 718 -924
rect 170 -994 172 -990
rect 499 -1018 501 -1008
rect 514 -1018 516 -1008
rect 534 -1018 536 -1008
rect 544 -1018 546 -1008
rect 570 -1018 572 -1008
rect 172 -1060 174 -1056
rect 358 -1093 360 -1083
rect 373 -1093 375 -1083
rect 393 -1093 395 -1083
rect 417 -1093 419 -1083
rect 175 -1127 177 -1123
rect 260 -1167 262 -1162
rect 281 -1167 283 -1162
rect 307 -1166 309 -1162
rect 175 -1194 177 -1190
<< ndiffusion >>
rect 407 -76 416 -70
rect 411 -80 416 -76
rect 418 -80 431 -70
rect 433 -80 446 -70
rect 448 -80 461 -70
rect 463 -80 475 -70
rect 477 -76 486 -70
rect 477 -80 482 -76
rect 492 -76 501 -70
rect 496 -80 501 -76
rect 503 -74 508 -70
rect 503 -80 512 -74
rect 169 -123 170 -119
rect 172 -123 173 -119
rect 857 -121 865 -118
rect 861 -125 865 -121
rect 867 -122 870 -118
rect 874 -122 877 -118
rect 867 -125 877 -122
rect 879 -121 892 -118
rect 879 -125 883 -121
rect 887 -125 892 -121
rect 894 -122 896 -118
rect 900 -122 902 -118
rect 894 -125 902 -122
rect 904 -122 909 -118
rect 904 -125 913 -122
rect 921 -122 925 -118
rect 917 -125 925 -122
rect 927 -122 930 -118
rect 927 -125 934 -122
rect 538 -176 547 -170
rect 542 -180 547 -176
rect 549 -180 562 -170
rect 564 -180 582 -170
rect 584 -180 592 -170
rect 594 -176 604 -170
rect 594 -180 600 -176
rect 609 -176 618 -170
rect 613 -180 618 -176
rect 620 -174 625 -170
rect 620 -180 629 -174
rect 171 -189 172 -185
rect 174 -189 175 -185
rect 174 -256 175 -252
rect 177 -256 178 -252
rect 174 -323 175 -319
rect 177 -323 178 -319
rect 192 -428 193 -424
rect 195 -428 196 -424
rect 88 -468 93 -467
rect 92 -472 93 -468
rect 95 -468 99 -467
rect 107 -468 112 -467
rect 95 -472 97 -468
rect 111 -472 112 -468
rect 114 -468 120 -467
rect 114 -472 116 -468
rect 132 -468 137 -467
rect 136 -472 137 -468
rect 139 -468 145 -467
rect 139 -472 141 -468
rect 151 -468 156 -467
rect 155 -472 156 -468
rect 158 -468 164 -467
rect 158 -472 160 -468
rect 194 -589 195 -585
rect 197 -589 198 -585
rect 90 -629 95 -628
rect 94 -633 95 -629
rect 97 -629 101 -628
rect 109 -629 114 -628
rect 97 -633 99 -629
rect 113 -633 114 -629
rect 116 -629 122 -628
rect 116 -633 118 -629
rect 134 -629 139 -628
rect 138 -633 139 -629
rect 141 -629 147 -628
rect 141 -633 143 -629
rect 153 -629 158 -628
rect 157 -633 158 -629
rect 160 -629 166 -628
rect 160 -633 162 -629
rect 676 -214 685 -208
rect 680 -218 685 -214
rect 687 -218 700 -208
rect 702 -218 720 -208
rect 722 -214 730 -208
rect 722 -218 726 -214
rect 735 -214 744 -208
rect 739 -218 744 -214
rect 746 -212 751 -208
rect 746 -218 755 -212
rect 857 -246 858 -242
rect 860 -246 861 -242
rect 809 -250 811 -246
rect 805 -253 811 -250
rect 813 -253 832 -246
rect 834 -249 841 -246
rect 834 -253 837 -249
rect 785 -650 794 -644
rect 789 -654 794 -650
rect 796 -654 809 -644
rect 811 -654 829 -644
rect 831 -654 839 -644
rect 841 -650 851 -644
rect 841 -654 847 -650
rect 856 -650 865 -644
rect 860 -654 865 -650
rect 867 -648 872 -644
rect 867 -654 876 -648
rect 193 -743 194 -739
rect 196 -743 197 -739
rect 89 -783 94 -782
rect 93 -787 94 -783
rect 96 -783 100 -782
rect 108 -783 113 -782
rect 96 -787 98 -783
rect 112 -787 113 -783
rect 115 -783 121 -782
rect 115 -787 117 -783
rect 133 -783 138 -782
rect 137 -787 138 -783
rect 140 -783 146 -782
rect 140 -787 142 -783
rect 152 -783 157 -782
rect 156 -787 157 -783
rect 159 -783 165 -782
rect 159 -787 161 -783
rect 193 -891 194 -887
rect 196 -891 197 -887
rect 848 -901 856 -898
rect 852 -905 856 -901
rect 858 -902 861 -898
rect 865 -902 868 -898
rect 858 -905 868 -902
rect 870 -901 883 -898
rect 870 -905 874 -901
rect 878 -905 883 -901
rect 885 -902 887 -898
rect 891 -902 893 -898
rect 885 -905 893 -902
rect 895 -902 900 -898
rect 895 -905 904 -902
rect 912 -902 916 -898
rect 908 -905 916 -902
rect 918 -902 921 -898
rect 918 -905 925 -902
rect 89 -931 94 -930
rect 93 -935 94 -931
rect 96 -931 100 -930
rect 108 -931 113 -930
rect 96 -935 98 -931
rect 112 -935 113 -931
rect 115 -931 121 -930
rect 115 -935 117 -931
rect 133 -931 138 -930
rect 137 -935 138 -931
rect 140 -931 146 -930
rect 140 -935 142 -931
rect 152 -931 157 -930
rect 156 -935 157 -931
rect 159 -931 165 -930
rect 159 -935 161 -931
rect 622 -965 631 -959
rect 626 -969 631 -965
rect 633 -969 646 -959
rect 648 -969 661 -959
rect 663 -969 676 -959
rect 678 -969 690 -959
rect 692 -965 701 -959
rect 692 -969 697 -965
rect 707 -965 716 -959
rect 711 -969 716 -965
rect 718 -963 723 -959
rect 718 -969 727 -963
rect 169 -1018 170 -1014
rect 172 -1018 173 -1014
rect 490 -1049 499 -1043
rect 494 -1053 499 -1049
rect 501 -1053 514 -1043
rect 516 -1053 534 -1043
rect 536 -1053 544 -1043
rect 546 -1049 556 -1043
rect 546 -1053 552 -1049
rect 561 -1049 570 -1043
rect 565 -1053 570 -1049
rect 572 -1047 577 -1043
rect 572 -1053 581 -1047
rect 171 -1084 172 -1080
rect 174 -1084 175 -1080
rect 349 -1124 358 -1118
rect 353 -1128 358 -1124
rect 360 -1128 373 -1118
rect 375 -1128 393 -1118
rect 395 -1124 403 -1118
rect 395 -1128 399 -1124
rect 408 -1124 417 -1118
rect 412 -1128 417 -1124
rect 419 -1122 424 -1118
rect 419 -1128 428 -1122
rect 174 -1151 175 -1147
rect 177 -1151 178 -1147
rect 306 -1190 307 -1186
rect 309 -1190 310 -1186
rect 258 -1194 260 -1190
rect 254 -1197 260 -1194
rect 262 -1197 281 -1190
rect 283 -1193 290 -1190
rect 283 -1197 286 -1193
rect 174 -1218 175 -1214
rect 177 -1218 178 -1214
<< pdiffusion >>
rect 407 -41 416 -35
rect 411 -45 416 -41
rect 418 -41 431 -35
rect 418 -45 420 -41
rect 424 -45 431 -41
rect 433 -41 446 -35
rect 433 -45 437 -41
rect 441 -45 446 -41
rect 448 -41 461 -35
rect 448 -45 452 -41
rect 456 -45 461 -41
rect 463 -41 475 -35
rect 463 -45 467 -41
rect 471 -45 475 -41
rect 477 -41 486 -35
rect 477 -45 482 -41
rect 492 -41 501 -35
rect 496 -45 501 -41
rect 503 -41 512 -35
rect 503 -45 508 -41
rect 169 -99 170 -95
rect 172 -99 173 -95
rect 538 -141 547 -135
rect 542 -145 547 -141
rect 549 -141 562 -135
rect 549 -145 553 -141
rect 558 -145 562 -141
rect 564 -141 582 -135
rect 564 -145 571 -141
rect 575 -145 582 -141
rect 584 -141 592 -135
rect 584 -145 586 -141
rect 590 -145 592 -141
rect 594 -141 604 -135
rect 594 -145 600 -141
rect 609 -141 618 -135
rect 613 -145 618 -141
rect 620 -141 629 -135
rect 620 -145 625 -141
rect 857 -91 865 -88
rect 861 -95 865 -91
rect 867 -95 877 -88
rect 879 -95 892 -88
rect 894 -95 902 -88
rect 904 -91 913 -88
rect 904 -95 909 -91
rect 917 -91 925 -88
rect 921 -95 925 -91
rect 927 -91 934 -88
rect 927 -95 930 -91
rect 171 -165 172 -161
rect 174 -165 175 -161
rect 676 -179 685 -173
rect 174 -232 175 -228
rect 177 -232 178 -228
rect 174 -299 175 -295
rect 177 -299 178 -295
rect 192 -404 193 -400
rect 195 -404 196 -400
rect 88 -437 93 -436
rect 92 -441 93 -437
rect 95 -437 101 -436
rect 95 -441 97 -437
rect 107 -437 112 -436
rect 111 -441 112 -437
rect 114 -437 120 -436
rect 114 -441 116 -437
rect 132 -437 137 -436
rect 136 -441 137 -437
rect 139 -437 145 -436
rect 139 -441 141 -437
rect 151 -437 156 -436
rect 155 -441 156 -437
rect 158 -437 164 -436
rect 158 -441 160 -437
rect 194 -565 195 -561
rect 197 -565 198 -561
rect 90 -598 95 -597
rect 94 -602 95 -598
rect 97 -598 103 -597
rect 97 -602 99 -598
rect 109 -598 114 -597
rect 113 -602 114 -598
rect 116 -598 122 -597
rect 116 -602 118 -598
rect 134 -598 139 -597
rect 138 -602 139 -598
rect 141 -598 147 -597
rect 141 -602 143 -598
rect 153 -598 158 -597
rect 157 -602 158 -598
rect 160 -598 166 -597
rect 160 -602 162 -598
rect 680 -183 685 -179
rect 687 -179 700 -173
rect 687 -183 691 -179
rect 696 -183 700 -179
rect 702 -179 720 -173
rect 702 -183 709 -179
rect 713 -183 720 -179
rect 722 -179 730 -173
rect 722 -183 726 -179
rect 735 -179 744 -173
rect 739 -183 744 -179
rect 746 -179 755 -173
rect 746 -183 751 -179
rect 805 -219 811 -218
rect 809 -223 811 -219
rect 813 -222 816 -218
rect 813 -223 820 -222
rect 826 -219 832 -218
rect 830 -223 832 -219
rect 834 -222 837 -218
rect 857 -222 858 -218
rect 860 -222 861 -218
rect 834 -223 841 -222
rect 785 -615 794 -609
rect 789 -619 794 -615
rect 796 -615 809 -609
rect 796 -619 800 -615
rect 805 -619 809 -615
rect 811 -615 829 -609
rect 811 -619 818 -615
rect 822 -619 829 -615
rect 831 -615 839 -609
rect 831 -619 833 -615
rect 837 -619 839 -615
rect 841 -615 851 -609
rect 841 -619 847 -615
rect 856 -615 865 -609
rect 860 -619 865 -615
rect 867 -615 876 -609
rect 867 -619 872 -615
rect 193 -719 194 -715
rect 196 -719 197 -715
rect 89 -752 94 -751
rect 93 -756 94 -752
rect 96 -752 102 -751
rect 96 -756 98 -752
rect 108 -752 113 -751
rect 112 -756 113 -752
rect 115 -752 121 -751
rect 115 -756 117 -752
rect 133 -752 138 -751
rect 137 -756 138 -752
rect 140 -752 146 -751
rect 140 -756 142 -752
rect 152 -752 157 -751
rect 156 -756 157 -752
rect 159 -752 165 -751
rect 159 -756 161 -752
rect 193 -867 194 -863
rect 196 -867 197 -863
rect 848 -871 856 -868
rect 852 -875 856 -871
rect 858 -875 868 -868
rect 870 -875 883 -868
rect 885 -875 893 -868
rect 895 -871 904 -868
rect 895 -875 900 -871
rect 908 -871 916 -868
rect 912 -875 916 -871
rect 918 -871 925 -868
rect 918 -875 921 -871
rect 89 -900 94 -899
rect 93 -904 94 -900
rect 96 -900 102 -899
rect 96 -904 98 -900
rect 108 -900 113 -899
rect 112 -904 113 -900
rect 115 -900 121 -899
rect 115 -904 117 -900
rect 133 -900 138 -899
rect 137 -904 138 -900
rect 140 -900 146 -899
rect 140 -904 142 -900
rect 152 -900 157 -899
rect 156 -904 157 -900
rect 159 -900 165 -899
rect 159 -904 161 -900
rect 622 -930 631 -924
rect 626 -934 631 -930
rect 633 -930 646 -924
rect 633 -934 635 -930
rect 639 -934 646 -930
rect 648 -930 661 -924
rect 648 -934 652 -930
rect 656 -934 661 -930
rect 663 -930 676 -924
rect 663 -934 667 -930
rect 671 -934 676 -930
rect 678 -930 690 -924
rect 678 -934 682 -930
rect 686 -934 690 -930
rect 692 -930 701 -924
rect 692 -934 697 -930
rect 707 -930 716 -924
rect 711 -934 716 -930
rect 718 -930 727 -924
rect 718 -934 723 -930
rect 169 -994 170 -990
rect 172 -994 173 -990
rect 490 -1014 499 -1008
rect 494 -1018 499 -1014
rect 501 -1014 514 -1008
rect 501 -1018 505 -1014
rect 510 -1018 514 -1014
rect 516 -1014 534 -1008
rect 516 -1018 523 -1014
rect 527 -1018 534 -1014
rect 536 -1014 544 -1008
rect 536 -1018 538 -1014
rect 542 -1018 544 -1014
rect 546 -1014 556 -1008
rect 546 -1018 552 -1014
rect 561 -1014 570 -1008
rect 565 -1018 570 -1014
rect 572 -1014 581 -1008
rect 572 -1018 577 -1014
rect 171 -1060 172 -1056
rect 174 -1060 175 -1056
rect 349 -1089 358 -1083
rect 353 -1093 358 -1089
rect 360 -1089 373 -1083
rect 360 -1093 364 -1089
rect 369 -1093 373 -1089
rect 375 -1089 393 -1083
rect 375 -1093 382 -1089
rect 386 -1093 393 -1089
rect 395 -1089 403 -1083
rect 395 -1093 399 -1089
rect 408 -1089 417 -1083
rect 412 -1093 417 -1089
rect 419 -1089 428 -1083
rect 419 -1093 424 -1089
rect 174 -1127 175 -1123
rect 177 -1127 178 -1123
rect 254 -1163 260 -1162
rect 258 -1167 260 -1163
rect 262 -1166 265 -1162
rect 262 -1167 269 -1166
rect 275 -1163 281 -1162
rect 279 -1167 281 -1163
rect 283 -1166 286 -1162
rect 306 -1166 307 -1162
rect 309 -1166 310 -1162
rect 283 -1167 290 -1166
rect 174 -1194 175 -1190
rect 177 -1194 178 -1190
<< ndcontact >>
rect 407 -80 411 -76
rect 482 -80 486 -76
rect 492 -80 496 -76
rect 508 -74 512 -70
rect 165 -123 169 -119
rect 173 -123 177 -119
rect 857 -125 861 -121
rect 870 -122 874 -118
rect 883 -125 887 -121
rect 896 -122 900 -118
rect 909 -122 913 -118
rect 917 -122 921 -118
rect 930 -122 934 -118
rect 538 -180 542 -176
rect 600 -180 604 -176
rect 609 -180 613 -176
rect 625 -174 629 -170
rect 167 -189 171 -185
rect 175 -189 179 -185
rect 170 -256 174 -252
rect 178 -256 182 -252
rect 170 -323 174 -319
rect 178 -323 182 -319
rect 188 -428 192 -424
rect 196 -428 200 -424
rect 88 -472 92 -468
rect 97 -472 101 -468
rect 107 -472 111 -468
rect 116 -472 120 -468
rect 132 -472 136 -468
rect 141 -472 145 -468
rect 151 -472 155 -468
rect 160 -472 164 -468
rect 190 -589 194 -585
rect 198 -589 202 -585
rect 90 -633 94 -629
rect 99 -633 103 -629
rect 109 -633 113 -629
rect 118 -633 122 -629
rect 134 -633 138 -629
rect 143 -633 147 -629
rect 153 -633 157 -629
rect 162 -633 166 -629
rect 676 -218 680 -214
rect 726 -218 730 -214
rect 735 -218 739 -214
rect 751 -212 755 -208
rect 853 -246 857 -242
rect 861 -246 865 -242
rect 805 -250 809 -246
rect 837 -253 841 -249
rect 785 -654 789 -650
rect 847 -654 851 -650
rect 856 -654 860 -650
rect 872 -648 876 -644
rect 189 -743 193 -739
rect 197 -743 201 -739
rect 89 -787 93 -783
rect 98 -787 102 -783
rect 108 -787 112 -783
rect 117 -787 121 -783
rect 133 -787 137 -783
rect 142 -787 146 -783
rect 152 -787 156 -783
rect 161 -787 165 -783
rect 189 -891 193 -887
rect 197 -891 201 -887
rect 848 -905 852 -901
rect 861 -902 865 -898
rect 874 -905 878 -901
rect 887 -902 891 -898
rect 900 -902 904 -898
rect 908 -902 912 -898
rect 921 -902 925 -898
rect 89 -935 93 -931
rect 98 -935 102 -931
rect 108 -935 112 -931
rect 117 -935 121 -931
rect 133 -935 137 -931
rect 142 -935 146 -931
rect 152 -935 156 -931
rect 161 -935 165 -931
rect 622 -969 626 -965
rect 697 -969 701 -965
rect 707 -969 711 -965
rect 723 -963 727 -959
rect 165 -1018 169 -1014
rect 173 -1018 177 -1014
rect 490 -1053 494 -1049
rect 552 -1053 556 -1049
rect 561 -1053 565 -1049
rect 577 -1047 581 -1043
rect 167 -1084 171 -1080
rect 175 -1084 179 -1080
rect 349 -1128 353 -1124
rect 399 -1128 403 -1124
rect 408 -1128 412 -1124
rect 424 -1122 428 -1118
rect 170 -1151 174 -1147
rect 178 -1151 182 -1147
rect 302 -1190 306 -1186
rect 310 -1190 314 -1186
rect 254 -1194 258 -1190
rect 286 -1197 290 -1193
rect 170 -1218 174 -1214
rect 178 -1218 182 -1214
<< pdcontact >>
rect 407 -45 411 -41
rect 420 -45 424 -41
rect 437 -45 441 -41
rect 452 -45 456 -41
rect 467 -45 471 -41
rect 482 -45 486 -41
rect 492 -45 496 -41
rect 508 -45 512 -41
rect 165 -99 169 -95
rect 173 -99 177 -95
rect 538 -145 542 -141
rect 553 -145 558 -141
rect 571 -145 575 -141
rect 586 -145 590 -141
rect 600 -145 604 -141
rect 609 -145 613 -141
rect 625 -145 629 -141
rect 857 -95 861 -91
rect 909 -95 913 -91
rect 917 -95 921 -91
rect 930 -95 934 -91
rect 167 -165 171 -161
rect 175 -165 179 -161
rect 170 -232 174 -228
rect 178 -232 182 -228
rect 170 -299 174 -295
rect 178 -299 182 -295
rect 188 -404 192 -400
rect 196 -404 200 -400
rect 88 -441 92 -437
rect 97 -441 101 -437
rect 107 -441 111 -437
rect 116 -441 120 -437
rect 132 -441 136 -437
rect 141 -441 145 -437
rect 151 -441 155 -437
rect 160 -441 164 -437
rect 190 -565 194 -561
rect 198 -565 202 -561
rect 90 -602 94 -598
rect 99 -602 103 -598
rect 109 -602 113 -598
rect 118 -602 122 -598
rect 134 -602 138 -598
rect 143 -602 147 -598
rect 153 -602 157 -598
rect 162 -602 166 -598
rect 676 -183 680 -179
rect 691 -183 696 -179
rect 709 -183 713 -179
rect 726 -183 730 -179
rect 735 -183 739 -179
rect 751 -183 755 -179
rect 805 -223 809 -219
rect 816 -222 820 -218
rect 826 -223 830 -219
rect 837 -222 841 -218
rect 853 -222 857 -218
rect 861 -222 865 -218
rect 785 -619 789 -615
rect 800 -619 805 -615
rect 818 -619 822 -615
rect 833 -619 837 -615
rect 847 -619 851 -615
rect 856 -619 860 -615
rect 872 -619 876 -615
rect 189 -719 193 -715
rect 197 -719 201 -715
rect 89 -756 93 -752
rect 98 -756 102 -752
rect 108 -756 112 -752
rect 117 -756 121 -752
rect 133 -756 137 -752
rect 142 -756 146 -752
rect 152 -756 156 -752
rect 161 -756 165 -752
rect 189 -867 193 -863
rect 197 -867 201 -863
rect 848 -875 852 -871
rect 900 -875 904 -871
rect 908 -875 912 -871
rect 921 -875 925 -871
rect 89 -904 93 -900
rect 98 -904 102 -900
rect 108 -904 112 -900
rect 117 -904 121 -900
rect 133 -904 137 -900
rect 142 -904 146 -900
rect 152 -904 156 -900
rect 161 -904 165 -900
rect 622 -934 626 -930
rect 635 -934 639 -930
rect 652 -934 656 -930
rect 667 -934 671 -930
rect 682 -934 686 -930
rect 697 -934 701 -930
rect 707 -934 711 -930
rect 723 -934 727 -930
rect 165 -994 169 -990
rect 173 -994 177 -990
rect 490 -1018 494 -1014
rect 505 -1018 510 -1014
rect 523 -1018 527 -1014
rect 538 -1018 542 -1014
rect 552 -1018 556 -1014
rect 561 -1018 565 -1014
rect 577 -1018 581 -1014
rect 167 -1060 171 -1056
rect 175 -1060 179 -1056
rect 349 -1093 353 -1089
rect 364 -1093 369 -1089
rect 382 -1093 386 -1089
rect 399 -1093 403 -1089
rect 408 -1093 412 -1089
rect 424 -1093 428 -1089
rect 170 -1127 174 -1123
rect 178 -1127 182 -1123
rect 254 -1167 258 -1163
rect 265 -1166 269 -1162
rect 275 -1167 279 -1163
rect 286 -1166 290 -1162
rect 302 -1166 306 -1162
rect 310 -1166 314 -1162
rect 170 -1194 174 -1190
rect 178 -1194 182 -1190
<< polysilicon >>
rect 416 -35 418 -32
rect 431 -35 433 -32
rect 446 -35 448 -32
rect 461 -35 463 -32
rect 475 -35 477 -32
rect 501 -35 503 -32
rect 416 -70 418 -45
rect 431 -70 433 -45
rect 446 -70 448 -45
rect 461 -70 463 -45
rect 475 -70 477 -45
rect 501 -61 503 -45
rect 518 -65 758 -61
rect 501 -70 503 -65
rect 170 -95 172 -92
rect 170 -112 172 -99
rect 416 -111 418 -80
rect 431 -99 433 -80
rect 446 -99 448 -80
rect 461 -99 463 -80
rect 475 -99 477 -80
rect 501 -83 503 -80
rect 34 -114 172 -112
rect 34 -946 36 -114
rect 170 -119 172 -114
rect 182 -115 418 -111
rect 170 -126 172 -123
rect 547 -135 549 -132
rect 562 -135 564 -132
rect 582 -135 584 -132
rect 592 -135 594 -132
rect 618 -135 620 -132
rect 755 -143 758 -65
rect 865 -88 867 -85
rect 877 -88 879 -85
rect 892 -88 894 -85
rect 902 -88 904 -85
rect 925 -88 927 -85
rect 865 -118 867 -95
rect 877 -118 879 -95
rect 892 -118 894 -95
rect 902 -118 904 -95
rect 925 -110 927 -95
rect 925 -118 927 -114
rect 865 -143 867 -125
rect 172 -161 174 -158
rect 172 -178 174 -165
rect 547 -170 549 -145
rect 562 -170 564 -145
rect 582 -170 584 -145
rect 592 -170 594 -145
rect 618 -161 620 -145
rect 755 -146 867 -143
rect 877 -161 879 -125
rect 635 -165 879 -161
rect 618 -170 620 -165
rect 41 -180 174 -178
rect 41 -798 43 -180
rect 172 -185 174 -180
rect 192 -181 517 -177
rect 685 -173 687 -170
rect 700 -173 702 -170
rect 720 -173 722 -170
rect 744 -173 746 -170
rect 172 -192 174 -189
rect 515 -199 517 -181
rect 547 -199 549 -180
rect 515 -201 549 -199
rect 175 -228 177 -225
rect 175 -245 177 -232
rect 48 -247 177 -245
rect 48 -644 50 -247
rect 175 -252 177 -247
rect 175 -259 177 -256
rect 175 -295 177 -292
rect 175 -312 177 -299
rect 65 -314 177 -312
rect 65 -483 67 -314
rect 175 -319 177 -314
rect 175 -326 177 -323
rect 193 -400 195 -397
rect 78 -407 114 -405
rect 65 -486 70 -483
rect 78 -492 80 -407
rect 93 -436 95 -433
rect 112 -436 114 -407
rect 193 -417 195 -404
rect 188 -419 195 -417
rect 193 -424 195 -419
rect 193 -431 195 -428
rect 137 -436 139 -433
rect 156 -436 158 -433
rect 93 -453 95 -441
rect 112 -444 114 -441
rect 137 -453 139 -441
rect 93 -455 114 -453
rect 93 -467 95 -464
rect 112 -467 114 -455
rect 138 -457 139 -453
rect 137 -467 139 -457
rect 156 -467 158 -441
rect 167 -456 173 -454
rect 93 -492 95 -472
rect 112 -483 114 -472
rect 137 -475 139 -472
rect 156 -483 158 -472
rect 116 -485 158 -483
rect 171 -492 173 -456
rect 78 -494 173 -492
rect 195 -561 197 -558
rect 80 -568 116 -566
rect 48 -647 72 -644
rect 80 -653 82 -568
rect 95 -597 97 -594
rect 114 -597 116 -568
rect 195 -578 197 -565
rect 190 -580 197 -578
rect 195 -585 197 -580
rect 195 -592 197 -589
rect 139 -597 141 -594
rect 158 -597 160 -594
rect 95 -614 97 -602
rect 114 -605 116 -602
rect 139 -614 141 -602
rect 95 -616 116 -614
rect 95 -628 97 -625
rect 114 -628 116 -616
rect 140 -618 141 -614
rect 139 -628 141 -618
rect 158 -628 160 -602
rect 169 -617 175 -615
rect 95 -653 97 -633
rect 114 -644 116 -633
rect 139 -636 141 -633
rect 158 -644 160 -633
rect 118 -646 160 -644
rect 173 -653 175 -617
rect 80 -655 175 -653
rect 562 -692 564 -180
rect 582 -199 584 -180
rect 592 -200 594 -180
rect 618 -183 620 -180
rect 685 -208 687 -183
rect 700 -208 702 -183
rect 720 -208 722 -183
rect 744 -199 746 -183
rect 892 -199 894 -125
rect 761 -203 894 -199
rect 744 -208 746 -203
rect 811 -218 813 -215
rect 832 -218 834 -215
rect 858 -218 860 -215
rect 685 -237 687 -218
rect 700 -259 702 -218
rect 720 -238 722 -218
rect 744 -221 746 -218
rect 811 -246 813 -223
rect 832 -246 834 -223
rect 858 -235 860 -222
rect 902 -234 904 -125
rect 925 -128 927 -125
rect 853 -237 860 -235
rect 858 -242 860 -237
rect 869 -238 904 -234
rect 858 -249 860 -246
rect 811 -311 813 -253
rect 832 -264 834 -253
rect 625 -315 813 -311
rect 794 -609 796 -606
rect 809 -609 811 -606
rect 829 -609 831 -606
rect 839 -609 841 -606
rect 865 -609 867 -606
rect 794 -644 796 -619
rect 809 -644 811 -619
rect 829 -644 831 -619
rect 839 -644 841 -619
rect 865 -635 867 -619
rect 865 -644 867 -639
rect 794 -671 796 -654
rect 771 -673 796 -671
rect 809 -678 811 -654
rect 771 -680 811 -678
rect 829 -686 831 -654
rect 771 -688 831 -686
rect 109 -696 564 -692
rect 839 -694 841 -654
rect 865 -657 867 -654
rect 771 -696 841 -694
rect 194 -715 196 -712
rect 79 -722 115 -720
rect 41 -801 71 -798
rect 79 -807 81 -722
rect 94 -751 96 -748
rect 113 -751 115 -722
rect 194 -732 196 -719
rect 189 -734 196 -732
rect 194 -739 196 -734
rect 194 -746 196 -743
rect 138 -751 140 -748
rect 157 -751 159 -748
rect 94 -768 96 -756
rect 113 -759 115 -756
rect 138 -768 140 -756
rect 94 -770 115 -768
rect 94 -782 96 -779
rect 113 -782 115 -770
rect 139 -772 140 -768
rect 138 -782 140 -772
rect 157 -782 159 -756
rect 168 -771 174 -769
rect 94 -807 96 -787
rect 113 -798 115 -787
rect 138 -790 140 -787
rect 157 -798 159 -787
rect 117 -800 159 -798
rect 172 -807 174 -771
rect 79 -809 174 -807
rect 194 -863 196 -860
rect 79 -870 115 -868
rect 34 -949 71 -946
rect 79 -955 81 -870
rect 94 -899 96 -896
rect 113 -899 115 -870
rect 194 -880 196 -867
rect 856 -868 858 -865
rect 868 -868 870 -865
rect 883 -868 885 -865
rect 893 -868 895 -865
rect 916 -868 918 -865
rect 189 -882 196 -880
rect 194 -887 196 -882
rect 194 -894 196 -891
rect 138 -899 140 -896
rect 157 -899 159 -896
rect 856 -898 858 -875
rect 868 -898 870 -875
rect 883 -898 885 -875
rect 893 -898 895 -875
rect 916 -890 918 -875
rect 916 -898 918 -894
rect 94 -916 96 -904
rect 113 -907 115 -904
rect 138 -916 140 -904
rect 94 -918 115 -916
rect 94 -930 96 -927
rect 113 -930 115 -918
rect 139 -920 140 -916
rect 138 -930 140 -920
rect 157 -930 159 -904
rect 168 -919 174 -917
rect 94 -955 96 -935
rect 113 -946 115 -935
rect 138 -938 140 -935
rect 157 -946 159 -935
rect 117 -948 159 -946
rect 172 -955 174 -919
rect 631 -924 633 -921
rect 646 -924 648 -921
rect 661 -924 663 -921
rect 676 -924 678 -921
rect 690 -924 692 -921
rect 716 -924 718 -921
rect 79 -957 174 -955
rect 631 -959 633 -934
rect 646 -959 648 -934
rect 661 -959 663 -934
rect 676 -959 678 -934
rect 690 -959 692 -934
rect 716 -950 718 -934
rect 856 -950 858 -905
rect 733 -954 858 -950
rect 716 -959 718 -954
rect 170 -990 172 -987
rect 631 -989 633 -969
rect 646 -989 648 -969
rect 661 -989 663 -969
rect 676 -988 678 -969
rect 690 -988 692 -969
rect 716 -972 718 -969
rect 409 -992 633 -989
rect 170 -1007 172 -994
rect 409 -1006 414 -992
rect 152 -1009 172 -1007
rect 170 -1014 172 -1009
rect 236 -1010 414 -1006
rect 499 -1008 501 -1005
rect 514 -1008 516 -1005
rect 534 -1008 536 -1005
rect 544 -1008 546 -1005
rect 570 -1008 572 -1005
rect 170 -1021 172 -1018
rect 499 -1043 501 -1018
rect 514 -1043 516 -1018
rect 534 -1043 536 -1018
rect 544 -1043 546 -1018
rect 570 -1034 572 -1018
rect 868 -1034 870 -905
rect 883 -918 885 -905
rect 587 -1038 870 -1034
rect 570 -1043 572 -1038
rect 172 -1056 174 -1053
rect 172 -1073 174 -1060
rect 499 -1072 501 -1053
rect 514 -1072 516 -1053
rect 534 -1071 536 -1053
rect 544 -1071 546 -1053
rect 570 -1056 572 -1053
rect 152 -1075 174 -1073
rect 172 -1080 174 -1075
rect 193 -1075 501 -1072
rect 358 -1083 360 -1080
rect 373 -1083 375 -1080
rect 393 -1083 395 -1080
rect 417 -1083 419 -1080
rect 172 -1087 174 -1084
rect 358 -1118 360 -1093
rect 373 -1118 375 -1093
rect 393 -1118 395 -1093
rect 417 -1109 419 -1093
rect 417 -1118 419 -1113
rect 175 -1123 177 -1120
rect 175 -1140 177 -1127
rect 152 -1142 177 -1140
rect 175 -1147 177 -1142
rect 187 -1143 340 -1139
rect 337 -1149 340 -1143
rect 358 -1149 360 -1128
rect 373 -1147 375 -1128
rect 175 -1154 177 -1151
rect 337 -1152 360 -1149
rect 393 -1148 395 -1128
rect 417 -1131 419 -1128
rect 260 -1162 262 -1159
rect 281 -1162 283 -1159
rect 307 -1162 309 -1159
rect 175 -1190 177 -1187
rect 260 -1190 262 -1167
rect 281 -1190 283 -1167
rect 307 -1179 309 -1166
rect 893 -1178 895 -905
rect 916 -908 918 -905
rect 302 -1181 309 -1179
rect 307 -1186 309 -1181
rect 318 -1182 895 -1178
rect 175 -1207 177 -1194
rect 307 -1193 309 -1190
rect 260 -1206 262 -1197
rect 152 -1209 177 -1207
rect 175 -1214 177 -1209
rect 188 -1210 262 -1206
rect 281 -1210 283 -1197
rect 175 -1221 177 -1218
<< polycontact >>
rect 499 -65 503 -61
rect 514 -65 518 -61
rect 430 -103 434 -99
rect 445 -103 449 -99
rect 460 -103 464 -99
rect 474 -103 478 -99
rect 178 -115 182 -111
rect 923 -114 927 -110
rect 616 -165 620 -161
rect 631 -165 635 -161
rect 188 -181 192 -177
rect 70 -487 74 -483
rect 184 -420 188 -416
rect 134 -457 138 -453
rect 163 -457 167 -453
rect 112 -487 116 -483
rect 72 -648 76 -644
rect 186 -581 190 -577
rect 136 -618 140 -614
rect 165 -618 169 -614
rect 114 -648 118 -644
rect 581 -203 585 -199
rect 591 -204 595 -200
rect 742 -203 746 -199
rect 757 -203 761 -199
rect 684 -241 688 -237
rect 719 -242 723 -238
rect 849 -238 853 -234
rect 865 -238 869 -234
rect 699 -263 703 -259
rect 831 -268 835 -264
rect 621 -315 625 -311
rect 863 -639 867 -635
rect 767 -673 771 -669
rect 767 -681 771 -677
rect 767 -689 771 -685
rect 105 -696 109 -692
rect 767 -697 771 -693
rect 71 -802 75 -798
rect 185 -735 189 -731
rect 135 -772 139 -768
rect 164 -772 168 -768
rect 113 -802 117 -798
rect 71 -950 75 -946
rect 185 -883 189 -879
rect 914 -894 918 -890
rect 135 -920 139 -916
rect 164 -920 168 -916
rect 113 -950 117 -946
rect 714 -954 718 -950
rect 729 -954 733 -950
rect 148 -1010 152 -1006
rect 645 -993 649 -989
rect 660 -993 664 -989
rect 675 -992 679 -988
rect 689 -992 693 -988
rect 232 -1010 236 -1006
rect 882 -922 886 -918
rect 568 -1038 572 -1034
rect 583 -1038 587 -1034
rect 148 -1076 152 -1072
rect 189 -1076 193 -1072
rect 513 -1076 517 -1072
rect 533 -1075 537 -1071
rect 543 -1075 547 -1071
rect 415 -1113 419 -1109
rect 148 -1143 152 -1139
rect 183 -1143 187 -1139
rect 372 -1151 376 -1147
rect 392 -1152 396 -1148
rect 298 -1182 302 -1178
rect 314 -1182 318 -1178
rect 148 -1210 152 -1206
rect 184 -1210 188 -1206
rect 280 -1214 284 -1210
<< metal1 >>
rect 371 -31 535 -28
rect 159 -90 170 -86
rect 371 -86 374 -31
rect 407 -41 411 -31
rect 437 -41 441 -31
rect 467 -41 471 -31
rect 492 -41 496 -31
rect 420 -61 424 -45
rect 452 -61 456 -45
rect 482 -61 486 -45
rect 508 -61 512 -45
rect 420 -65 499 -61
rect 508 -65 514 -61
rect 482 -76 486 -65
rect 508 -70 512 -65
rect 175 -89 374 -86
rect 407 -86 411 -80
rect 492 -86 496 -80
rect 532 -80 535 -31
rect 532 -83 921 -80
rect 407 -89 523 -86
rect 175 -90 184 -89
rect 165 -95 168 -90
rect 173 -111 176 -99
rect 407 -101 411 -89
rect 208 -105 411 -101
rect 173 -115 178 -111
rect 173 -119 176 -115
rect 166 -128 169 -123
rect 208 -128 211 -105
rect 430 -106 434 -103
rect 445 -106 449 -103
rect 460 -106 464 -103
rect 474 -106 478 -103
rect 165 -131 178 -128
rect 183 -131 211 -128
rect 161 -156 169 -152
rect 174 -156 186 -152
rect 167 -161 170 -156
rect 175 -177 178 -165
rect 175 -181 188 -177
rect 175 -185 178 -181
rect 168 -194 171 -189
rect 520 -190 523 -89
rect 532 -128 535 -83
rect 857 -91 861 -83
rect 917 -91 921 -83
rect 909 -110 913 -95
rect 930 -106 934 -95
rect 930 -110 939 -106
rect 870 -114 923 -110
rect 870 -118 874 -114
rect 896 -118 900 -114
rect 930 -118 934 -110
rect 532 -131 653 -128
rect 538 -141 542 -131
rect 571 -141 575 -131
rect 600 -141 604 -131
rect 609 -141 613 -131
rect 553 -161 558 -145
rect 586 -161 590 -145
rect 625 -161 629 -145
rect 553 -165 616 -161
rect 625 -165 631 -161
rect 600 -176 604 -165
rect 625 -170 629 -165
rect 650 -166 653 -131
rect 857 -130 861 -125
rect 883 -130 887 -125
rect 909 -130 913 -122
rect 917 -130 921 -122
rect 857 -133 921 -130
rect 650 -169 783 -166
rect 538 -190 542 -180
rect 609 -190 613 -180
rect 676 -179 680 -169
rect 709 -179 713 -169
rect 735 -179 739 -169
rect 520 -193 650 -190
rect 167 -197 178 -194
rect 164 -223 169 -219
rect 174 -223 189 -219
rect 581 -216 585 -203
rect 449 -219 585 -216
rect 170 -228 173 -223
rect 591 -223 595 -204
rect 464 -226 595 -223
rect 647 -228 650 -193
rect 691 -199 696 -183
rect 726 -199 730 -183
rect 751 -199 755 -183
rect 691 -203 742 -199
rect 751 -203 757 -199
rect 726 -214 730 -203
rect 751 -208 755 -203
rect 780 -209 783 -169
rect 780 -213 872 -209
rect 676 -228 680 -218
rect 735 -228 739 -218
rect 805 -219 809 -213
rect 647 -231 773 -228
rect 178 -244 181 -232
rect 240 -241 684 -237
rect 240 -244 244 -241
rect 178 -248 244 -244
rect 178 -252 181 -248
rect 719 -250 723 -242
rect 450 -253 723 -250
rect 770 -256 773 -231
rect 816 -239 820 -222
rect 826 -219 830 -213
rect 853 -218 856 -213
rect 837 -239 841 -222
rect 861 -234 864 -222
rect 844 -238 849 -234
rect 861 -238 865 -234
rect 844 -239 847 -238
rect 816 -243 847 -239
rect 861 -242 864 -238
rect 805 -256 809 -250
rect 837 -249 841 -243
rect 854 -256 857 -246
rect 914 -256 917 -133
rect 171 -261 174 -256
rect 770 -259 917 -256
rect 170 -264 178 -261
rect 164 -290 169 -286
rect 174 -290 189 -286
rect 170 -295 173 -290
rect 178 -311 181 -299
rect 178 -315 621 -311
rect 178 -319 181 -315
rect 171 -328 174 -323
rect 170 -331 178 -328
rect 151 -395 169 -391
rect 88 -413 128 -409
rect 88 -437 92 -413
rect 88 -454 92 -441
rect 75 -457 92 -454
rect 88 -468 92 -457
rect 97 -420 116 -416
rect 97 -437 101 -420
rect 116 -437 120 -421
rect 97 -468 101 -441
rect 107 -468 111 -441
rect 116 -468 120 -441
rect 124 -453 128 -413
rect 151 -421 155 -395
rect 174 -395 207 -391
rect 188 -400 191 -395
rect 196 -416 199 -404
rect 182 -420 184 -416
rect 196 -420 306 -416
rect 132 -425 155 -421
rect 196 -424 199 -420
rect 132 -437 136 -425
rect 151 -437 155 -425
rect 189 -433 192 -428
rect 177 -436 192 -433
rect 124 -457 134 -453
rect 141 -461 145 -441
rect 124 -465 145 -461
rect 107 -475 111 -472
rect 124 -475 128 -465
rect 141 -468 145 -465
rect 160 -453 164 -441
rect 160 -457 163 -453
rect 160 -468 164 -457
rect 107 -479 128 -475
rect 132 -475 136 -472
rect 151 -475 155 -472
rect 177 -474 182 -436
rect 177 -475 178 -474
rect 132 -479 178 -475
rect 74 -486 112 -483
rect 74 -496 77 -486
rect 20 -499 77 -496
rect 20 -1243 23 -499
rect 153 -556 169 -552
rect 90 -574 130 -570
rect 90 -598 94 -574
rect 90 -615 94 -602
rect 77 -618 94 -615
rect 90 -629 94 -618
rect 99 -581 118 -577
rect 99 -598 103 -581
rect 118 -598 122 -582
rect 99 -629 103 -602
rect 109 -629 113 -602
rect 118 -629 122 -602
rect 126 -614 130 -574
rect 153 -582 157 -556
rect 174 -556 204 -552
rect 190 -561 193 -556
rect 198 -577 201 -565
rect 184 -581 186 -577
rect 198 -579 268 -577
rect 134 -586 157 -582
rect 198 -582 269 -579
rect 198 -585 201 -582
rect 134 -598 138 -586
rect 153 -598 157 -586
rect 191 -594 194 -589
rect 126 -618 136 -614
rect 143 -622 147 -602
rect 126 -626 147 -622
rect 109 -636 113 -633
rect 126 -636 130 -626
rect 143 -629 147 -626
rect 162 -614 166 -602
rect 184 -597 194 -594
rect 162 -618 165 -614
rect 162 -629 166 -618
rect 109 -640 130 -636
rect 134 -636 138 -633
rect 153 -636 157 -633
rect 179 -636 184 -599
rect 134 -640 184 -636
rect 76 -647 114 -644
rect 76 -654 79 -647
rect 260 -648 269 -582
rect 297 -628 306 -420
rect 699 -527 703 -263
rect 831 -275 835 -268
rect 351 -530 703 -527
rect 782 -605 882 -602
rect 785 -615 789 -605
rect 818 -615 822 -605
rect 847 -615 851 -605
rect 856 -615 860 -605
rect 297 -633 444 -628
rect 449 -633 743 -628
rect 298 -634 743 -633
rect 38 -657 79 -654
rect 260 -653 459 -648
rect 464 -653 722 -648
rect 260 -655 722 -653
rect 260 -656 269 -655
rect 38 -1100 41 -657
rect 719 -677 722 -655
rect 740 -670 743 -634
rect 800 -635 805 -619
rect 833 -635 837 -619
rect 872 -635 876 -619
rect 800 -639 863 -635
rect 872 -639 881 -635
rect 847 -650 851 -639
rect 872 -644 876 -639
rect 785 -664 789 -654
rect 856 -664 860 -654
rect 785 -667 855 -664
rect 740 -673 767 -670
rect 719 -680 767 -677
rect 621 -688 767 -685
rect 94 -696 105 -692
rect 152 -710 169 -706
rect 89 -728 129 -724
rect 89 -752 93 -728
rect 89 -769 93 -756
rect 76 -772 93 -769
rect 89 -783 93 -772
rect 98 -735 117 -731
rect 98 -752 102 -735
rect 117 -752 121 -736
rect 98 -783 102 -756
rect 108 -783 112 -756
rect 117 -783 121 -756
rect 125 -768 129 -728
rect 152 -736 156 -710
rect 174 -710 208 -706
rect 189 -715 192 -710
rect 197 -731 200 -719
rect 183 -735 185 -731
rect 197 -735 473 -731
rect 621 -731 624 -688
rect 478 -735 624 -731
rect 693 -697 767 -694
rect 133 -740 156 -736
rect 197 -739 200 -735
rect 133 -752 137 -740
rect 152 -752 156 -740
rect 190 -748 193 -743
rect 125 -772 135 -768
rect 142 -776 146 -756
rect 125 -780 146 -776
rect 108 -790 112 -787
rect 125 -790 129 -780
rect 142 -783 146 -780
rect 161 -768 165 -756
rect 183 -751 193 -748
rect 161 -772 164 -768
rect 161 -783 165 -772
rect 108 -794 129 -790
rect 133 -790 137 -787
rect 152 -790 156 -787
rect 178 -790 183 -753
rect 133 -794 183 -790
rect 75 -801 113 -798
rect 75 -809 78 -801
rect 49 -812 78 -809
rect 49 -1036 52 -812
rect 152 -858 169 -854
rect 89 -876 129 -872
rect 89 -900 93 -876
rect 89 -917 93 -904
rect 76 -920 93 -917
rect 89 -931 93 -920
rect 98 -883 117 -879
rect 98 -900 102 -883
rect 117 -900 121 -884
rect 98 -931 102 -904
rect 108 -931 112 -904
rect 117 -931 121 -904
rect 125 -916 129 -876
rect 152 -884 156 -858
rect 174 -858 208 -854
rect 189 -863 192 -858
rect 197 -879 200 -867
rect 693 -879 699 -697
rect 183 -883 185 -879
rect 197 -883 699 -879
rect 789 -863 912 -860
rect 133 -888 156 -884
rect 197 -887 200 -883
rect 133 -900 137 -888
rect 152 -900 156 -888
rect 190 -896 193 -891
rect 125 -920 135 -916
rect 142 -924 146 -904
rect 125 -928 146 -924
rect 108 -938 112 -935
rect 125 -938 129 -928
rect 142 -931 146 -928
rect 161 -916 165 -904
rect 183 -899 193 -896
rect 161 -920 164 -916
rect 161 -931 165 -920
rect 108 -942 129 -938
rect 133 -938 137 -935
rect 152 -938 156 -935
rect 178 -938 183 -901
rect 789 -917 792 -863
rect 848 -871 852 -863
rect 908 -871 912 -863
rect 900 -890 904 -875
rect 921 -886 925 -875
rect 921 -890 930 -886
rect 861 -894 914 -890
rect 861 -898 865 -894
rect 887 -898 891 -894
rect 921 -898 925 -890
rect 848 -910 852 -905
rect 874 -910 878 -905
rect 900 -910 904 -902
rect 908 -910 912 -902
rect 848 -913 912 -910
rect 618 -920 792 -917
rect 622 -930 626 -920
rect 652 -930 656 -920
rect 682 -930 686 -920
rect 707 -930 711 -920
rect 133 -942 183 -938
rect 75 -949 113 -946
rect 75 -963 78 -949
rect 635 -950 639 -934
rect 667 -950 671 -934
rect 697 -950 701 -934
rect 723 -950 727 -934
rect 635 -954 714 -950
rect 723 -954 729 -950
rect 75 -966 617 -963
rect 697 -965 701 -954
rect 723 -959 727 -954
rect 159 -985 169 -981
rect 174 -985 184 -981
rect 165 -990 168 -985
rect 173 -1006 176 -994
rect 584 -1001 587 -980
rect 612 -996 617 -966
rect 622 -975 626 -969
rect 707 -975 711 -969
rect 861 -975 864 -913
rect 882 -928 886 -922
rect 622 -978 864 -975
rect 645 -996 649 -993
rect 612 -999 649 -996
rect 487 -1004 587 -1001
rect 129 -1010 148 -1006
rect 173 -1010 232 -1006
rect 173 -1014 176 -1010
rect 490 -1014 494 -1004
rect 523 -1014 527 -1004
rect 552 -1014 556 -1004
rect 561 -1014 565 -1004
rect 166 -1023 169 -1018
rect 165 -1026 178 -1023
rect 505 -1034 510 -1018
rect 538 -1034 542 -1018
rect 577 -1034 581 -1018
rect 49 -1040 472 -1036
rect 505 -1038 568 -1034
rect 577 -1038 583 -1034
rect 161 -1051 169 -1047
rect 174 -1051 186 -1047
rect 167 -1056 170 -1051
rect 175 -1072 178 -1060
rect 129 -1076 148 -1072
rect 175 -1076 189 -1072
rect 175 -1080 178 -1076
rect 346 -1079 430 -1076
rect 168 -1089 171 -1084
rect 349 -1089 353 -1079
rect 382 -1089 386 -1079
rect 408 -1089 412 -1079
rect 468 -1080 472 -1040
rect 552 -1049 556 -1038
rect 577 -1043 581 -1038
rect 490 -1063 494 -1053
rect 561 -1063 565 -1053
rect 652 -1063 655 -978
rect 660 -1001 664 -993
rect 490 -1066 655 -1063
rect 513 -1080 517 -1076
rect 468 -1083 517 -1080
rect 523 -1088 527 -1066
rect 533 -1081 537 -1075
rect 543 -1081 547 -1075
rect 167 -1092 178 -1089
rect 38 -1103 337 -1100
rect 164 -1118 169 -1114
rect 174 -1118 189 -1114
rect 170 -1123 173 -1118
rect 178 -1139 181 -1127
rect 121 -1143 148 -1139
rect 178 -1143 183 -1139
rect 178 -1147 181 -1143
rect 171 -1156 174 -1151
rect 170 -1159 178 -1156
rect 233 -1157 317 -1153
rect 164 -1185 169 -1181
rect 233 -1181 236 -1157
rect 254 -1163 258 -1157
rect 174 -1185 236 -1181
rect 265 -1183 269 -1166
rect 275 -1163 279 -1157
rect 302 -1162 305 -1157
rect 334 -1157 337 -1103
rect 364 -1109 369 -1093
rect 399 -1109 403 -1093
rect 424 -1109 428 -1093
rect 478 -1091 527 -1088
rect 364 -1113 415 -1109
rect 424 -1113 431 -1109
rect 399 -1124 403 -1113
rect 424 -1118 428 -1113
rect 349 -1138 353 -1128
rect 408 -1138 412 -1128
rect 478 -1138 481 -1091
rect 518 -1102 521 -1100
rect 675 -1102 679 -992
rect 689 -1000 693 -992
rect 518 -1105 679 -1102
rect 349 -1141 481 -1138
rect 372 -1157 376 -1151
rect 334 -1160 376 -1157
rect 286 -1183 290 -1166
rect 310 -1178 313 -1166
rect 293 -1182 298 -1178
rect 310 -1182 314 -1178
rect 293 -1183 296 -1182
rect 170 -1190 173 -1185
rect 265 -1187 296 -1183
rect 310 -1186 313 -1182
rect 178 -1206 181 -1194
rect 254 -1201 258 -1194
rect 286 -1193 290 -1187
rect 303 -1201 306 -1190
rect 383 -1201 386 -1141
rect 392 -1156 396 -1152
rect 254 -1204 386 -1201
rect 100 -1210 148 -1206
rect 178 -1210 184 -1206
rect 178 -1214 181 -1210
rect 171 -1223 174 -1218
rect 269 -1223 272 -1204
rect 170 -1226 178 -1223
rect 183 -1226 272 -1223
rect 280 -1243 284 -1214
rect 20 -1246 284 -1243
<< m2contact >>
rect 429 -111 434 -106
rect 444 -111 449 -106
rect 459 -111 464 -106
rect 473 -111 478 -106
rect 444 -220 449 -215
rect 459 -227 464 -222
rect 445 -254 450 -249
rect 70 -459 75 -454
rect 116 -421 121 -416
rect 177 -420 182 -415
rect 72 -620 77 -615
rect 118 -582 123 -577
rect 179 -581 184 -576
rect 346 -532 351 -527
rect 444 -633 449 -628
rect 459 -653 464 -648
rect 89 -697 94 -692
rect 71 -774 76 -769
rect 117 -736 122 -731
rect 178 -735 183 -730
rect 473 -735 478 -730
rect 71 -922 76 -917
rect 117 -884 122 -879
rect 178 -883 183 -878
rect 613 -922 618 -917
rect 583 -980 588 -975
rect 124 -1010 129 -1005
rect 124 -1077 129 -1072
rect 341 -1081 346 -1076
rect 659 -1006 664 -1001
rect 532 -1086 537 -1081
rect 542 -1086 547 -1081
rect 116 -1144 121 -1139
rect 317 -1158 322 -1153
rect 516 -1100 521 -1095
rect 688 -1005 693 -1000
rect 392 -1161 397 -1156
rect 95 -1211 100 -1206
<< metal2 >>
rect 430 -116 434 -111
rect 445 -116 449 -111
rect 460 -113 464 -111
rect 474 -113 478 -111
rect 54 -376 372 -373
rect 54 -454 59 -376
rect 121 -420 177 -416
rect 182 -420 183 -416
rect 27 -457 70 -454
rect 27 -1206 30 -457
rect 56 -530 346 -527
rect 56 -615 59 -530
rect 123 -581 179 -577
rect 184 -581 185 -577
rect 44 -618 72 -615
rect 44 -1139 47 -618
rect 54 -696 89 -692
rect 54 -769 57 -696
rect 122 -735 178 -731
rect 183 -735 184 -731
rect 54 -772 71 -769
rect 54 -1072 57 -772
rect 430 -844 433 -116
rect 445 -215 448 -116
rect 445 -249 448 -220
rect 460 -222 463 -113
rect 445 -628 448 -254
rect 62 -847 433 -844
rect 62 -917 65 -847
rect 122 -883 178 -879
rect 183 -883 184 -879
rect 62 -920 71 -917
rect 62 -1006 65 -920
rect 62 -1010 124 -1006
rect 54 -1076 124 -1072
rect 317 -1079 341 -1076
rect 44 -1143 116 -1139
rect 317 -1153 321 -1079
rect 445 -1139 448 -633
rect 460 -648 463 -227
rect 460 -1095 463 -653
rect 474 -730 477 -113
rect 474 -990 477 -735
rect 584 -920 613 -917
rect 584 -975 587 -920
rect 474 -993 615 -990
rect 612 -1001 615 -993
rect 612 -1004 659 -1001
rect 533 -1095 537 -1086
rect 460 -1098 516 -1095
rect 521 -1098 537 -1095
rect 543 -1139 547 -1086
rect 689 -1139 693 -1005
rect 445 -1142 693 -1139
rect 445 -1156 448 -1142
rect 397 -1159 448 -1156
rect 27 -1210 95 -1206
<< m3contact >>
rect 372 -378 377 -373
<< m123contact >>
rect 170 -90 175 -85
rect 178 -133 183 -128
rect 169 -156 174 -151
rect 178 -199 183 -194
rect 169 -223 174 -218
rect 178 -266 183 -261
rect 169 -290 174 -285
rect 178 -333 183 -328
rect 169 -396 174 -391
rect 178 -479 183 -474
rect 169 -557 174 -552
rect 204 -557 209 -552
rect 179 -599 184 -594
rect 169 -711 174 -706
rect 178 -753 183 -748
rect 169 -859 174 -854
rect 178 -901 183 -896
rect 169 -985 174 -980
rect 178 -1028 183 -1023
rect 169 -1051 174 -1046
rect 178 -1094 183 -1089
rect 169 -1118 174 -1113
rect 430 -1081 435 -1076
rect 431 -1114 436 -1109
rect 830 -280 835 -275
rect 777 -607 782 -602
rect 855 -669 860 -664
rect 881 -933 886 -928
rect 482 -1006 487 -1001
rect 178 -1161 183 -1156
rect 169 -1185 174 -1180
rect 178 -1228 183 -1223
<< metal3 >>
rect 170 -151 174 -90
rect 170 -218 174 -156
rect 170 -285 174 -223
rect 170 -391 174 -290
rect 170 -552 174 -396
rect 170 -706 174 -557
rect 170 -854 174 -711
rect 170 -980 174 -859
rect 170 -1046 174 -985
rect 170 -1113 174 -1051
rect 170 -1180 174 -1118
rect 178 -194 182 -133
rect 178 -261 182 -199
rect 178 -328 182 -266
rect 178 -474 182 -333
rect 831 -373 835 -280
rect 377 -377 835 -373
rect 178 -594 182 -479
rect 209 -556 777 -552
rect 178 -599 179 -594
rect 178 -748 182 -599
rect 773 -605 777 -556
rect 178 -766 182 -753
rect 856 -766 860 -669
rect 178 -769 860 -766
rect 178 -896 182 -769
rect 178 -1023 182 -901
rect 431 -1004 482 -1001
rect 178 -1089 182 -1028
rect 431 -1076 434 -1004
rect 178 -1156 182 -1094
rect 882 -1109 886 -933
rect 436 -1113 886 -1109
rect 178 -1223 182 -1161
<< labels >>
rlabel metal1 75 -455 75 -455 1 a3
rlabel metal1 77 -616 77 -616 1 a2
rlabel metal1 77 -645 77 -645 1 b2
rlabel metal1 76 -770 76 -770 1 a1
rlabel metal1 75 -799 75 -799 1 b1
rlabel metal1 76 -919 76 -919 1 a0
rlabel metal1 76 -948 76 -948 1 b0
rlabel metal1 74 -485 74 -485 1 b3
rlabel metal1 183 -313 183 -313 1 b3n
rlabel metal1 184 -246 184 -246 1 b2n
rlabel metal1 178 -113 178 -113 1 b0n
rlabel metal1 180 -179 180 -179 1 b1n
rlabel metal1 177 -1008 177 -1008 1 a0n
rlabel metal1 177 -1074 177 -1074 1 a1n
rlabel polycontact 184 -1141 184 -1141 1 a2n
rlabel metal1 184 -1208 184 -1208 1 a3n
rlabel metal1 937 -108 937 -108 7 gtr
rlabel metal1 155 -709 155 -709 1 VDD
rlabel metal1 164 -793 164 -793 1 gnd
rlabel metal1 879 -637 879 -637 1 equ
rlabel metal1 928 -888 928 -888 1 lsr
rlabel polysilicon 857 -916 857 -916 1 w1
rlabel polysilicon 869 -916 869 -916 1 w2
rlabel polysilicon 884 -916 884 -916 1 w3
rlabel polysilicon 894 -916 894 -916 1 w4
<< end >>
