magic
tech scmos
timestamp 1700230136
<< nwell >>
rect 2919 664 3021 685
rect 3114 665 3216 686
rect 3327 664 3429 685
rect 3528 665 3630 686
<< ntransistor >>
rect 2930 640 2932 645
rect 2956 640 2958 645
rect 2981 640 2983 645
rect 3007 640 3009 645
rect 3125 641 3127 646
rect 3151 641 3153 646
rect 3176 641 3178 646
rect 3202 641 3204 646
rect 3338 640 3340 645
rect 3364 640 3366 645
rect 3389 640 3391 645
rect 3415 640 3417 645
rect 3539 641 3541 646
rect 3565 641 3567 646
rect 3590 641 3592 646
rect 3616 641 3618 646
<< ptransistor >>
rect 2930 671 2932 676
rect 2956 671 2958 676
rect 2981 671 2983 676
rect 3007 671 3009 676
rect 3125 672 3127 677
rect 3151 672 3153 677
rect 3176 672 3178 677
rect 3202 672 3204 677
rect 3338 671 3340 676
rect 3364 671 3366 676
rect 3389 671 3391 676
rect 3415 671 3417 676
rect 3539 672 3541 677
rect 3565 672 3567 677
rect 3590 672 3592 677
rect 3616 672 3618 677
<< ndiffusion >>
rect 2929 641 2930 645
rect 2925 640 2930 641
rect 2932 641 2934 645
rect 2932 640 2938 641
rect 2955 641 2956 645
rect 2951 640 2956 641
rect 2958 641 2960 645
rect 2958 640 2964 641
rect 2976 644 2981 645
rect 2980 640 2981 644
rect 2983 641 2986 645
rect 2983 640 2990 641
rect 3001 644 3007 645
rect 3005 640 3007 644
rect 3009 641 3010 645
rect 3009 640 3014 641
rect 3124 642 3125 646
rect 3120 641 3125 642
rect 3127 642 3129 646
rect 3127 641 3133 642
rect 3150 642 3151 646
rect 3146 641 3151 642
rect 3153 642 3155 646
rect 3153 641 3159 642
rect 3171 645 3176 646
rect 3175 641 3176 645
rect 3178 642 3181 646
rect 3178 641 3185 642
rect 3196 645 3202 646
rect 3200 641 3202 645
rect 3204 642 3205 646
rect 3204 641 3209 642
rect 3337 641 3338 645
rect 3333 640 3338 641
rect 3340 641 3342 645
rect 3340 640 3346 641
rect 3363 641 3364 645
rect 3359 640 3364 641
rect 3366 641 3368 645
rect 3366 640 3372 641
rect 3384 644 3389 645
rect 3388 640 3389 644
rect 3391 641 3394 645
rect 3391 640 3398 641
rect 3409 644 3415 645
rect 3413 640 3415 644
rect 3417 641 3418 645
rect 3417 640 3422 641
rect 3538 642 3539 646
rect 3534 641 3539 642
rect 3541 642 3543 646
rect 3541 641 3547 642
rect 3564 642 3565 646
rect 3560 641 3565 642
rect 3567 642 3569 646
rect 3567 641 3573 642
rect 3585 645 3590 646
rect 3589 641 3590 645
rect 3592 642 3595 646
rect 3592 641 3599 642
rect 3610 645 3616 646
rect 3614 641 3616 645
rect 3618 642 3619 646
rect 3618 641 3623 642
<< pdiffusion >>
rect 2925 675 2930 676
rect 2929 671 2930 675
rect 2932 675 2938 676
rect 2932 671 2934 675
rect 2951 675 2956 676
rect 2955 671 2956 675
rect 2958 675 2964 676
rect 2958 671 2960 675
rect 2980 672 2981 676
rect 2976 671 2981 672
rect 2983 675 2990 676
rect 2983 671 2986 675
rect 3005 673 3007 676
rect 3001 671 3007 673
rect 3009 675 3014 676
rect 3009 671 3010 675
rect 3120 676 3125 677
rect 3124 672 3125 676
rect 3127 676 3133 677
rect 3127 672 3129 676
rect 3146 676 3151 677
rect 3150 672 3151 676
rect 3153 676 3159 677
rect 3153 672 3155 676
rect 3175 673 3176 677
rect 3171 672 3176 673
rect 3178 676 3185 677
rect 3178 672 3181 676
rect 3200 674 3202 677
rect 3196 672 3202 674
rect 3204 676 3209 677
rect 3204 672 3205 676
rect 3333 675 3338 676
rect 3337 671 3338 675
rect 3340 675 3346 676
rect 3340 671 3342 675
rect 3359 675 3364 676
rect 3363 671 3364 675
rect 3366 675 3372 676
rect 3366 671 3368 675
rect 3388 672 3389 676
rect 3384 671 3389 672
rect 3391 675 3398 676
rect 3391 671 3394 675
rect 3413 673 3415 676
rect 3409 671 3415 673
rect 3417 675 3422 676
rect 3417 671 3418 675
rect 3534 676 3539 677
rect 3538 672 3539 676
rect 3541 676 3547 677
rect 3541 672 3543 676
rect 3560 676 3565 677
rect 3564 672 3565 676
rect 3567 676 3573 677
rect 3567 672 3569 676
rect 3589 673 3590 677
rect 3585 672 3590 673
rect 3592 676 3599 677
rect 3592 672 3595 676
rect 3614 674 3616 677
rect 3610 672 3616 674
rect 3618 676 3623 677
rect 3618 672 3619 676
<< ndcontact >>
rect 2925 641 2929 645
rect 2934 641 2938 645
rect 2951 641 2955 645
rect 2960 641 2964 645
rect 2976 640 2980 644
rect 2986 641 2990 645
rect 3001 640 3005 644
rect 3010 641 3014 645
rect 3120 642 3124 646
rect 3129 642 3133 646
rect 3146 642 3150 646
rect 3155 642 3159 646
rect 3171 641 3175 645
rect 3181 642 3185 646
rect 3196 641 3200 645
rect 3205 642 3209 646
rect 3333 641 3337 645
rect 3342 641 3346 645
rect 3359 641 3363 645
rect 3368 641 3372 645
rect 3384 640 3388 644
rect 3394 641 3398 645
rect 3409 640 3413 644
rect 3418 641 3422 645
rect 3534 642 3538 646
rect 3543 642 3547 646
rect 3560 642 3564 646
rect 3569 642 3573 646
rect 3585 641 3589 645
rect 3595 642 3599 646
rect 3610 641 3614 645
rect 3619 642 3623 646
<< pdcontact >>
rect 2925 671 2929 675
rect 2934 671 2938 675
rect 2951 671 2955 675
rect 2960 671 2964 675
rect 2976 672 2980 676
rect 2986 671 2990 675
rect 3001 673 3005 677
rect 3010 671 3014 675
rect 3120 672 3124 676
rect 3129 672 3133 676
rect 3146 672 3150 676
rect 3155 672 3159 676
rect 3171 673 3175 677
rect 3181 672 3185 676
rect 3196 674 3200 678
rect 3205 672 3209 676
rect 3333 671 3337 675
rect 3342 671 3346 675
rect 3359 671 3363 675
rect 3368 671 3372 675
rect 3384 672 3388 676
rect 3394 671 3398 675
rect 3409 673 3413 677
rect 3418 671 3422 675
rect 3534 672 3538 676
rect 3543 672 3547 676
rect 3560 672 3564 676
rect 3569 672 3573 676
rect 3585 673 3589 677
rect 3595 672 3599 676
rect 3610 674 3614 678
rect 3619 672 3623 676
<< polysilicon >>
rect 2807 713 2988 717
rect 3007 717 3009 721
rect 3099 717 3183 718
rect 2993 714 3183 717
rect 2993 713 3098 714
rect 3202 718 3204 722
rect 3188 717 3322 718
rect 3415 717 3417 721
rect 3530 717 3597 718
rect 3188 714 3396 717
rect 2915 686 2958 688
rect 2859 583 2864 656
rect 2915 630 2917 686
rect 2930 676 2932 681
rect 2956 676 2958 686
rect 2981 676 2983 679
rect 3007 676 3009 713
rect 3110 687 3153 689
rect 2930 662 2932 671
rect 2956 668 2958 671
rect 2930 660 2958 662
rect 2930 645 2932 648
rect 2956 645 2958 660
rect 2981 659 2983 671
rect 2981 645 2983 655
rect 3007 645 3009 671
rect 3017 657 3023 659
rect 2930 630 2932 640
rect 2915 628 2932 630
rect 2930 624 2932 628
rect 2956 629 2958 640
rect 2981 637 2983 640
rect 3007 629 3009 640
rect 2956 627 3009 629
rect 3021 624 3023 657
rect 3110 631 3112 687
rect 3125 677 3127 682
rect 3151 677 3153 687
rect 3176 677 3178 682
rect 3202 677 3204 714
rect 3312 713 3396 714
rect 3401 714 3597 717
rect 3401 713 3532 714
rect 3323 686 3366 688
rect 3125 663 3127 672
rect 3151 669 3153 672
rect 3125 661 3153 663
rect 3125 646 3127 649
rect 3151 646 3153 661
rect 3176 660 3178 672
rect 3176 646 3178 656
rect 3202 646 3204 672
rect 3212 658 3218 660
rect 3125 631 3127 641
rect 3110 629 3127 631
rect 2930 622 3023 624
rect 3125 625 3127 629
rect 3151 630 3153 641
rect 3176 638 3178 641
rect 3202 630 3204 641
rect 3151 628 3204 630
rect 3216 625 3218 658
rect 3125 623 3218 625
rect 3305 593 3308 636
rect 3323 630 3325 686
rect 3338 676 3340 681
rect 3364 676 3366 686
rect 3389 676 3391 680
rect 3415 676 3417 713
rect 3338 662 3340 671
rect 3364 668 3366 671
rect 3338 660 3366 662
rect 3338 645 3340 648
rect 3364 645 3366 660
rect 3389 659 3391 671
rect 3389 645 3391 655
rect 3415 645 3417 671
rect 3425 657 3431 659
rect 3338 630 3340 640
rect 3323 628 3340 630
rect 3338 624 3340 628
rect 3364 629 3366 640
rect 3389 637 3391 640
rect 3415 629 3417 640
rect 3364 627 3417 629
rect 3429 624 3431 657
rect 3338 622 3431 624
rect 3512 583 3517 700
rect 3524 687 3567 689
rect 3524 631 3526 687
rect 3539 677 3541 682
rect 3565 677 3567 687
rect 3590 677 3592 680
rect 3616 677 3618 722
rect 3539 663 3541 672
rect 3565 669 3567 672
rect 3539 661 3567 663
rect 3539 646 3541 649
rect 3565 646 3567 661
rect 3590 660 3592 672
rect 3590 646 3592 656
rect 3616 646 3618 672
rect 3626 658 3632 660
rect 3539 631 3541 641
rect 3524 629 3541 631
rect 3539 625 3541 629
rect 3565 630 3567 641
rect 3590 638 3592 641
rect 3616 630 3618 641
rect 3565 628 3618 630
rect 3630 625 3632 658
rect 3539 623 3632 625
rect 2859 577 3517 583
<< polycontact >>
rect 3005 721 3011 727
rect 3200 722 3206 728
rect 2988 712 2993 718
rect 3183 713 3188 719
rect 3413 721 3419 727
rect 3614 722 3620 728
rect 2857 656 2865 663
rect 2979 655 2983 659
rect 3013 656 3017 660
rect 3396 712 3401 717
rect 3597 713 3602 719
rect 3174 656 3178 660
rect 3208 657 3212 661
rect 3303 636 3310 643
rect 3510 700 3517 706
rect 3387 655 3391 659
rect 3421 656 3425 660
rect 3304 587 3310 593
rect 3588 656 3592 660
rect 3622 657 3626 661
<< metal1 >>
rect 3198 727 3200 728
rect 3003 726 3005 727
rect 2849 721 2885 726
rect 2892 721 3005 726
rect 3011 723 3200 727
rect 3099 722 3200 723
rect 3612 727 3614 728
rect 3411 726 3413 727
rect 3206 722 3413 726
rect 3312 721 3413 722
rect 3419 722 3614 727
rect 2849 708 2853 721
rect 3396 717 3401 718
rect 2861 708 2867 709
rect 2861 704 2929 708
rect 2861 703 2867 704
rect 2925 700 2972 704
rect 2925 675 2929 700
rect 2823 658 2857 662
rect 2925 645 2929 671
rect 2934 692 2964 696
rect 2934 675 2938 692
rect 2960 675 2964 692
rect 2934 645 2938 671
rect 2951 645 2955 671
rect 2960 645 2964 671
rect 2968 659 2972 700
rect 2988 691 2991 712
rect 3098 707 3124 710
rect 3120 705 3124 707
rect 3120 701 3167 705
rect 2976 687 3005 691
rect 2976 676 2980 687
rect 3001 677 3005 687
rect 3120 676 3124 701
rect 2968 655 2979 659
rect 2986 651 2990 671
rect 2968 647 2990 651
rect 2951 638 2955 641
rect 2968 638 2972 647
rect 2986 645 2990 647
rect 2951 634 2972 638
rect 3010 660 3014 671
rect 3010 656 3013 660
rect 3010 645 3014 656
rect 2976 637 2980 640
rect 3120 646 3124 672
rect 3129 693 3159 697
rect 3129 676 3133 693
rect 3155 676 3159 693
rect 3129 646 3133 672
rect 3146 646 3150 672
rect 3155 646 3159 672
rect 3163 660 3167 701
rect 3183 692 3186 713
rect 3305 700 3380 704
rect 3171 688 3200 692
rect 3171 677 3175 688
rect 3196 678 3200 688
rect 3163 656 3174 660
rect 3181 652 3185 672
rect 3163 648 3185 652
rect 3001 637 3005 640
rect 2976 633 3005 637
rect 3146 639 3150 642
rect 3163 639 3167 648
rect 3181 646 3185 648
rect 3146 635 3167 639
rect 3205 661 3209 672
rect 3205 657 3208 661
rect 3205 646 3209 657
rect 3171 638 3175 641
rect 3305 643 3308 700
rect 3333 675 3337 700
rect 3333 645 3337 671
rect 3196 638 3200 641
rect 3171 634 3200 638
rect 3342 692 3372 696
rect 3342 675 3346 692
rect 3368 675 3372 692
rect 3342 645 3346 671
rect 3359 645 3363 671
rect 3368 645 3372 671
rect 3376 659 3380 700
rect 3396 691 3399 712
rect 3517 701 3581 705
rect 3384 687 3413 691
rect 3384 676 3388 687
rect 3409 677 3413 687
rect 3534 676 3538 701
rect 3376 655 3387 659
rect 3394 651 3398 671
rect 3376 647 3398 651
rect 3359 638 3363 641
rect 3376 638 3380 647
rect 3394 645 3398 647
rect 3359 634 3380 638
rect 3418 660 3422 671
rect 3418 656 3421 660
rect 3418 645 3422 656
rect 3384 637 3388 640
rect 3534 646 3538 672
rect 3543 693 3573 697
rect 3543 676 3547 693
rect 3569 676 3573 693
rect 3543 646 3547 672
rect 3560 646 3564 672
rect 3569 646 3573 672
rect 3577 660 3581 701
rect 3597 692 3600 713
rect 3585 688 3614 692
rect 3585 677 3589 688
rect 3610 678 3614 688
rect 3577 656 3588 660
rect 3595 652 3599 672
rect 3577 648 3599 652
rect 3409 637 3413 640
rect 2992 619 2996 633
rect 3187 619 3191 634
rect 3384 633 3413 637
rect 3560 639 3564 642
rect 3577 639 3581 648
rect 3595 646 3599 648
rect 3560 635 3581 639
rect 3619 661 3623 672
rect 3619 657 3622 661
rect 3619 646 3623 657
rect 3585 638 3589 641
rect 3610 638 3614 641
rect 3585 634 3614 638
rect 3400 619 3404 633
rect 3601 619 3605 634
rect 2992 618 3191 619
rect 3399 618 3605 619
rect 2818 615 3605 618
rect 2818 614 3105 615
rect 3312 614 3534 615
rect 2825 587 3304 591
<< m2contact >>
rect 3090 704 3098 711
<< metal2 >>
rect 3092 611 3096 704
rect 2862 607 3096 611
<< labels >>
rlabel metal1 2948 693 2948 694 1 gbu3
rlabel metal1 3143 694 3143 695 1 gbu2
rlabel metal1 3358 693 3358 694 1 gbu1
rlabel metal1 3556 694 3556 695 1 gbu0
<< end >>
