magic
tech scmos
timestamp 1698930151
<< nwell >>
rect 66 -15 168 6
<< ntransistor >>
rect 77 -39 79 -34
rect 103 -39 105 -34
rect 128 -39 130 -34
rect 154 -39 156 -34
<< ptransistor >>
rect 77 -8 79 -3
rect 103 -8 105 -3
rect 128 -8 130 -3
rect 154 -8 156 -3
<< ndiffusion >>
rect 76 -38 77 -34
rect 72 -39 77 -38
rect 79 -38 81 -34
rect 79 -39 85 -38
rect 102 -38 103 -34
rect 98 -39 103 -38
rect 105 -38 107 -34
rect 105 -39 111 -38
rect 123 -35 128 -34
rect 127 -39 128 -35
rect 130 -38 133 -34
rect 130 -39 137 -38
rect 148 -35 154 -34
rect 152 -39 154 -35
rect 156 -38 157 -34
rect 156 -39 161 -38
<< pdiffusion >>
rect 72 -4 77 -3
rect 76 -8 77 -4
rect 79 -4 85 -3
rect 79 -8 81 -4
rect 98 -4 103 -3
rect 102 -8 103 -4
rect 105 -4 111 -3
rect 105 -8 107 -4
rect 127 -7 128 -3
rect 123 -8 128 -7
rect 130 -4 137 -3
rect 130 -8 133 -4
rect 152 -6 154 -3
rect 148 -8 154 -6
rect 156 -4 161 -3
rect 156 -8 157 -4
<< ndcontact >>
rect 72 -38 76 -34
rect 81 -38 85 -34
rect 98 -38 102 -34
rect 107 -38 111 -34
rect 123 -39 127 -35
rect 133 -38 137 -34
rect 148 -39 152 -35
rect 157 -38 161 -34
<< pdcontact >>
rect 72 -8 76 -4
rect 81 -8 85 -4
rect 98 -8 102 -4
rect 107 -8 111 -4
rect 123 -7 127 -3
rect 133 -8 137 -4
rect 148 -6 152 -2
rect 157 -8 161 -4
<< polysilicon >>
rect 62 7 105 9
rect 62 -49 64 7
rect 77 -3 79 2
rect 103 -3 105 7
rect 128 -3 130 0
rect 154 -3 156 1
rect 77 -17 79 -8
rect 103 -11 105 -8
rect 77 -19 105 -17
rect 77 -34 79 -31
rect 103 -34 105 -19
rect 128 -20 130 -8
rect 128 -34 130 -24
rect 154 -34 156 -8
rect 164 -22 170 -20
rect 77 -49 79 -39
rect 62 -51 79 -49
rect 77 -55 79 -51
rect 103 -50 105 -39
rect 128 -42 130 -39
rect 154 -50 156 -39
rect 103 -52 156 -50
rect 168 -55 170 -22
rect 77 -57 170 -55
<< polycontact >>
rect 126 -24 130 -20
rect 160 -23 164 -19
<< metal1 >>
rect 72 21 119 25
rect 72 -4 76 21
rect 72 -34 76 -8
rect 81 13 111 17
rect 81 -4 85 13
rect 107 -4 111 13
rect 81 -34 85 -8
rect 98 -34 102 -8
rect 107 -34 111 -8
rect 115 -20 119 21
rect 123 8 152 12
rect 123 -3 127 8
rect 148 -2 152 8
rect 115 -24 126 -20
rect 133 -28 137 -8
rect 115 -32 137 -28
rect 98 -41 102 -38
rect 115 -41 119 -32
rect 133 -34 137 -32
rect 98 -45 119 -41
rect 157 -19 161 -8
rect 157 -23 160 -19
rect 157 -34 161 -23
rect 123 -42 127 -39
rect 148 -42 152 -39
rect 123 -46 152 -42
<< labels >>
rlabel polysilicon 129 -18 129 -18 1 A
rlabel polysilicon 155 -23 155 -23 1 B
rlabel metal1 137 -44 137 -44 1 gnd
rlabel metal1 136 9 136 9 1 vdd
rlabel metal1 90 15 90 15 1 out
<< end >>
