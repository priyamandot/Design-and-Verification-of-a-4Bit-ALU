magic
tech scmos
timestamp 1698914331
<< nwell >>
rect -332 242 -263 261
rect -254 242 -227 261
<< ntransistor >>
rect -321 218 -319 223
rect -312 218 -310 223
rect -303 218 -301 223
rect -294 218 -292 223
rect -285 218 -283 223
rect -243 218 -241 223
<< ptransistor >>
rect -321 249 -319 254
rect -312 249 -310 254
rect -303 249 -301 254
rect -294 249 -292 254
rect -285 249 -283 254
rect -243 249 -241 254
<< ndiffusion >>
rect -326 222 -321 223
rect -322 218 -321 222
rect -319 218 -312 223
rect -310 218 -303 223
rect -301 218 -294 223
rect -292 218 -285 223
rect -283 219 -281 223
rect -277 219 -269 223
rect -283 218 -269 219
rect -248 221 -243 223
rect -244 218 -243 221
rect -241 220 -238 223
rect -241 218 -234 220
<< pdiffusion >>
rect -322 251 -321 254
rect -326 249 -321 251
rect -319 252 -312 254
rect -319 249 -317 252
rect -313 249 -312 252
rect -310 251 -308 254
rect -304 251 -303 254
rect -310 249 -303 251
rect -301 252 -294 254
rect -301 249 -299 252
rect -295 249 -294 252
rect -292 251 -290 254
rect -286 251 -285 254
rect -292 249 -285 251
rect -283 252 -269 254
rect -283 249 -281 252
rect -277 249 -269 252
rect -244 251 -243 254
rect -248 249 -243 251
rect -241 250 -238 254
rect -241 249 -234 250
<< ndcontact >>
rect -326 218 -322 222
rect -281 219 -277 223
rect -248 217 -244 221
rect -238 220 -234 224
<< pdcontact >>
rect -326 251 -322 255
rect -317 248 -313 252
rect -308 251 -304 255
rect -299 248 -295 252
rect -290 251 -286 255
rect -281 248 -277 252
rect -248 251 -244 255
rect -238 250 -234 254
<< polysilicon >>
rect -321 254 -319 257
rect -312 254 -310 257
rect -321 223 -319 249
rect -303 254 -301 257
rect -294 254 -292 257
rect -312 223 -310 249
rect -303 223 -301 249
rect -285 254 -283 257
rect -294 223 -292 249
rect -285 223 -283 249
rect -243 254 -241 257
rect -243 238 -241 249
rect -242 234 -241 238
rect -243 223 -241 234
rect -321 215 -319 218
rect -312 215 -310 218
rect -303 215 -301 218
rect -294 215 -292 218
rect -285 215 -283 218
rect -243 215 -241 218
<< polycontact >>
rect -246 234 -242 238
<< metal1 >>
rect -331 258 -230 261
rect -326 255 -322 258
rect -308 255 -304 258
rect -290 255 -286 258
rect -317 238 -313 248
rect -248 255 -244 258
rect -299 238 -295 248
rect -281 238 -277 248
rect -238 238 -234 250
rect -317 234 -246 238
rect -238 234 -230 238
rect -281 223 -277 234
rect -238 224 -234 234
rect -326 214 -322 218
rect -248 214 -244 217
rect -331 211 -230 214
<< labels >>
rlabel metal1 -308 212 -308 212 1 gnd
rlabel metal1 -294 260 -294 260 5 vdd
rlabel polysilicon -320 235 -320 235 1 A
rlabel polysilicon -311 232 -311 232 1 B
rlabel polysilicon -302 232 -302 232 1 C
rlabel polysilicon -293 232 -293 232 1 D
rlabel polysilicon -284 232 -284 232 1 E
rlabel metal1 -230 234 -230 238 7 out
<< end >>
