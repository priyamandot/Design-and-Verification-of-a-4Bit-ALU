magic
tech scmos
timestamp 1700301932
<< nwell >>
rect 73 214 98 231
rect 3 139 105 160
<< ntransistor >>
rect 85 197 87 201
rect 14 115 16 120
rect 40 115 42 120
rect 65 115 67 120
rect 91 115 93 120
<< ptransistor >>
rect 85 220 87 224
rect 14 146 16 151
rect 40 146 42 151
rect 65 146 67 151
rect 91 146 93 151
<< ndiffusion >>
rect 84 197 85 201
rect 87 197 88 201
rect 13 116 14 120
rect 9 115 14 116
rect 16 116 18 120
rect 16 115 22 116
rect 39 116 40 120
rect 35 115 40 116
rect 42 116 44 120
rect 42 115 48 116
rect 60 119 65 120
rect 64 115 65 119
rect 67 116 70 120
rect 67 115 74 116
rect 85 119 91 120
rect 89 115 91 119
rect 93 116 94 120
rect 93 115 98 116
<< pdiffusion >>
rect 84 220 85 224
rect 87 220 88 224
rect 9 150 14 151
rect 13 146 14 150
rect 16 150 22 151
rect 16 146 18 150
rect 35 150 40 151
rect 39 146 40 150
rect 42 150 48 151
rect 42 146 44 150
rect 64 147 65 151
rect 60 146 65 147
rect 67 150 74 151
rect 67 146 70 150
rect 89 148 91 151
rect 85 146 91 148
rect 93 150 98 151
rect 93 146 94 150
<< ndcontact >>
rect 80 197 84 201
rect 88 197 92 201
rect 9 116 13 120
rect 18 116 22 120
rect 35 116 39 120
rect 44 116 48 120
rect 60 115 64 119
rect 70 116 74 120
rect 85 115 89 119
rect 94 116 98 120
<< pdcontact >>
rect 80 220 84 224
rect 88 220 92 224
rect 9 146 13 150
rect 18 146 22 150
rect 35 146 39 150
rect 44 146 48 150
rect 60 147 64 151
rect 70 146 74 150
rect 85 148 89 152
rect 94 146 98 150
<< polysilicon >>
rect 34 172 37 205
rect 66 166 69 228
rect 85 224 87 227
rect 85 210 87 220
rect 81 208 87 210
rect 85 201 87 208
rect 85 194 87 197
rect -1 161 42 163
rect -1 105 1 161
rect 14 151 16 156
rect 40 151 42 161
rect 65 151 67 154
rect 91 151 93 155
rect 14 137 16 146
rect 40 143 42 146
rect 14 135 42 137
rect 14 120 16 123
rect 40 120 42 135
rect 65 134 67 146
rect 65 120 67 130
rect 91 120 93 146
rect 101 132 107 134
rect 14 105 16 115
rect -1 103 16 105
rect 14 99 16 103
rect 40 104 42 115
rect 65 112 67 115
rect 91 104 93 115
rect 40 102 93 104
rect 105 99 107 132
rect 14 97 107 99
<< polycontact >>
rect 65 228 69 232
rect 33 205 39 212
rect 33 167 38 172
rect 77 207 81 211
rect 66 162 70 166
rect 63 130 67 134
rect 97 131 101 135
<< metal1 >>
rect 69 228 98 231
rect 81 224 84 228
rect 88 211 92 220
rect 39 207 77 211
rect 88 207 95 211
rect 88 201 92 207
rect 81 193 84 197
rect 74 190 122 193
rect 9 175 56 179
rect 9 150 13 175
rect 9 120 13 146
rect 18 167 33 171
rect 38 167 48 171
rect 18 150 22 167
rect 44 150 48 167
rect 18 120 22 146
rect 35 120 39 146
rect 44 120 48 146
rect 52 134 56 175
rect 60 162 66 166
rect 70 162 89 166
rect 60 151 64 162
rect 85 152 89 162
rect 52 130 63 134
rect 70 126 74 146
rect 52 122 74 126
rect 35 113 39 116
rect 52 113 56 122
rect 70 120 74 122
rect 35 109 56 113
rect 94 135 98 146
rect 94 131 97 135
rect 94 120 98 131
rect 60 112 64 115
rect 85 112 89 115
rect 60 108 89 112
rect 75 95 78 108
rect 119 95 122 190
rect 75 92 122 95
<< labels >>
rlabel polysilicon 66 136 66 136 1 A
rlabel polysilicon 92 131 92 131 1 B
rlabel metal1 74 110 74 110 1 gnd
rlabel metal1 73 163 73 163 1 vdd
rlabel metal1 95 207 95 211 1 xnor_out
<< end >>
