magic
tech scmos
timestamp 1700302380
<< nwell >>
rect 0 99 52 118
rect 61 99 88 118
<< ntransistor >>
rect 11 75 13 80
rect 20 75 22 80
rect 29 75 31 80
rect 72 75 74 80
<< ptransistor >>
rect 11 106 13 111
rect 20 106 22 111
rect 29 106 31 111
rect 72 106 74 111
<< ndiffusion >>
rect 6 79 11 80
rect 10 75 11 79
rect 13 75 20 80
rect 22 75 29 80
rect 31 79 38 80
rect 31 75 33 79
rect 37 75 38 79
rect 67 78 72 80
rect 71 75 72 78
rect 74 77 77 80
rect 74 75 81 77
<< pdiffusion >>
rect 10 108 11 111
rect 6 106 11 108
rect 13 109 20 111
rect 13 106 15 109
rect 19 106 20 109
rect 22 108 24 111
rect 28 108 29 111
rect 22 106 29 108
rect 31 109 38 111
rect 31 106 33 109
rect 37 106 38 109
rect 71 108 72 111
rect 67 106 72 108
rect 74 107 77 111
rect 74 106 81 107
<< ndcontact >>
rect 6 75 10 79
rect 33 75 37 79
rect 67 74 71 78
rect 77 77 81 81
<< pdcontact >>
rect 6 108 10 112
rect 15 105 19 109
rect 24 108 28 112
rect 33 105 37 109
rect 67 108 71 112
rect 77 107 81 111
<< polysilicon >>
rect 11 111 13 114
rect 20 111 22 114
rect 11 80 13 106
rect 29 111 31 114
rect 20 80 22 106
rect 29 80 31 106
rect 72 111 74 114
rect 72 95 74 106
rect 73 91 74 95
rect 72 80 74 91
rect 11 72 13 75
rect 20 72 22 75
rect 29 72 31 75
rect 72 72 74 75
<< polycontact >>
rect 69 91 73 95
<< metal1 >>
rect 1 115 85 118
rect 6 112 10 115
rect 24 112 28 115
rect 67 112 71 115
rect 15 95 19 105
rect 33 95 37 105
rect 77 95 81 107
rect 15 91 69 95
rect 77 91 85 95
rect 33 79 37 91
rect 77 81 81 91
rect 6 71 10 75
rect 67 71 71 74
rect 1 68 85 71
<< labels >>
rlabel metal1 24 69 24 69 1 gnd
rlabel polysilicon 12 92 12 92 1 A
rlabel polysilicon 21 89 21 89 1 B
rlabel polysilicon 30 89 30 89 1 C
rlabel metal1 85 91 85 95 7 out
rlabel metal1 58 117 58 117 5 vdd
<< end >>
