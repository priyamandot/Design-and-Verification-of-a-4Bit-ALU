magic
tech scmos
timestamp 1700331077
<< nwell >>
rect 202 3538 304 3559
rect 379 3539 481 3560
rect 765 3545 867 3566
rect 942 3546 1044 3567
rect 1962 3562 2064 3583
rect 2139 3563 2241 3584
rect 1341 3531 1443 3552
rect 1518 3532 1620 3553
rect 227 3447 263 3466
rect 270 3447 297 3466
rect 413 3453 449 3472
rect 456 3453 483 3472
rect 544 3460 591 3479
rect 600 3460 627 3479
rect 790 3454 826 3473
rect 833 3454 860 3473
rect 976 3460 1012 3479
rect 1019 3460 1046 3479
rect 1107 3467 1154 3486
rect 1163 3467 1190 3486
rect 1366 3440 1402 3459
rect 1409 3440 1436 3459
rect 1552 3446 1588 3465
rect 1595 3446 1622 3465
rect 1683 3453 1730 3472
rect 1739 3453 1766 3472
rect 1987 3471 2023 3490
rect 2030 3471 2057 3490
rect 2173 3477 2209 3496
rect 2216 3477 2243 3496
rect 2304 3484 2351 3503
rect 2360 3484 2387 3503
rect 2959 3238 3061 3259
rect 3136 3239 3238 3260
rect 3522 3245 3624 3266
rect 3699 3246 3801 3267
rect 4719 3262 4821 3283
rect 4896 3263 4998 3284
rect 4098 3231 4200 3252
rect 4275 3232 4377 3253
rect 2984 3147 3020 3166
rect 3027 3147 3054 3166
rect 3170 3153 3206 3172
rect 3213 3153 3240 3172
rect 3301 3160 3348 3179
rect 3357 3160 3384 3179
rect 3547 3154 3583 3173
rect 3590 3154 3617 3173
rect 3733 3160 3769 3179
rect 3776 3160 3803 3179
rect 3864 3167 3911 3186
rect 3920 3167 3947 3186
rect 4123 3140 4159 3159
rect 4166 3140 4193 3159
rect 4309 3146 4345 3165
rect 4352 3146 4379 3165
rect 4440 3153 4487 3172
rect 4496 3153 4523 3172
rect 4744 3171 4780 3190
rect 4787 3171 4814 3190
rect 4930 3177 4966 3196
rect 4973 3177 5000 3196
rect 5061 3184 5108 3203
rect 5117 3184 5144 3203
rect 386 3047 424 3066
rect 431 3047 458 3066
rect 529 3047 567 3066
rect 574 3047 601 3066
rect 692 3047 730 3066
rect 737 3047 764 3066
rect 848 3047 886 3066
rect 893 3047 920 3066
rect 986 3047 1024 3066
rect 1031 3047 1058 3066
rect 1129 3047 1167 3066
rect 1174 3047 1201 3066
rect 1292 3047 1330 3066
rect 1337 3047 1364 3066
rect 1448 3047 1486 3066
rect 1493 3047 1520 3066
rect 230 2979 266 2998
rect 273 2979 300 2998
rect 182 2928 207 2945
rect 1686 2928 1788 2949
rect 1881 2929 1983 2950
rect 2094 2928 2196 2949
rect 2295 2929 2397 2950
rect 94 2895 129 2914
rect 136 2895 163 2914
rect 227 2898 265 2917
rect 272 2898 299 2917
rect 386 2905 424 2924
rect 431 2905 458 2924
rect 529 2905 567 2924
rect 574 2905 601 2924
rect 692 2905 730 2924
rect 737 2905 764 2924
rect 848 2905 886 2924
rect 893 2905 920 2924
rect 986 2905 1024 2924
rect 1031 2905 1058 2924
rect 1129 2905 1167 2924
rect 1174 2905 1201 2924
rect 1292 2905 1330 2924
rect 1337 2905 1364 2924
rect 1448 2905 1486 2924
rect 1493 2905 1520 2924
rect 182 2845 207 2862
rect 231 2807 269 2826
rect 276 2807 303 2826
rect 386 2756 424 2775
rect 431 2756 458 2775
rect 529 2756 567 2775
rect 574 2756 601 2775
rect 692 2756 730 2775
rect 737 2756 764 2775
rect 848 2756 886 2775
rect 893 2756 920 2775
rect 986 2756 1024 2775
rect 1031 2756 1058 2775
rect 1129 2756 1167 2775
rect 1174 2756 1201 2775
rect 1292 2756 1330 2775
rect 1337 2756 1364 2775
rect 1448 2756 1486 2775
rect 1493 2756 1520 2775
rect 2354 2736 2471 2759
rect 2112 2682 2137 2701
rect 2804 2686 2893 2707
rect 386 2631 424 2650
rect 431 2631 458 2650
rect 529 2631 567 2650
rect 574 2631 601 2650
rect 692 2631 730 2650
rect 737 2631 764 2650
rect 848 2631 886 2650
rect 893 2631 920 2650
rect 986 2631 1024 2650
rect 1031 2631 1058 2650
rect 1129 2631 1167 2650
rect 1174 2631 1201 2650
rect 1292 2631 1330 2650
rect 1337 2631 1364 2650
rect 1448 2631 1486 2650
rect 1493 2631 1520 2650
rect 2485 2636 2588 2659
rect 2114 2616 2139 2635
rect 2623 2598 2714 2621
rect 2117 2549 2142 2568
rect 2752 2557 2825 2578
rect 2117 2482 2142 2501
rect 2135 2377 2160 2396
rect 2034 2337 2125 2360
rect 768 2272 806 2291
rect 813 2272 840 2291
rect 911 2272 949 2291
rect 956 2272 983 2291
rect 1074 2272 1112 2291
rect 1119 2272 1146 2291
rect 1230 2272 1268 2291
rect 1275 2272 1302 2291
rect 2137 2216 2162 2235
rect 2036 2176 2127 2199
rect 2732 2162 2835 2185
rect 2895 2157 2931 2176
rect 2937 2157 2964 2176
rect 2136 2062 2161 2081
rect 2035 2022 2126 2045
rect 2136 1914 2161 1933
rect 2795 1906 2884 1927
rect 2035 1874 2126 1897
rect 2569 1847 2686 1870
rect 2112 1787 2137 1806
rect 2437 1763 2540 1786
rect 2114 1721 2139 1740
rect 2296 1688 2387 1711
rect 2117 1654 2142 1673
rect 2201 1613 2274 1634
rect 2117 1587 2142 1606
<< ntransistor >>
rect 213 3514 215 3519
rect 239 3514 241 3519
rect 264 3514 266 3519
rect 290 3514 292 3519
rect 390 3515 392 3520
rect 416 3515 418 3520
rect 441 3515 443 3520
rect 467 3515 469 3520
rect 776 3521 778 3526
rect 802 3521 804 3526
rect 827 3521 829 3526
rect 853 3521 855 3526
rect 953 3522 955 3527
rect 979 3522 981 3527
rect 1004 3522 1006 3527
rect 1030 3522 1032 3527
rect 1352 3507 1354 3512
rect 1378 3507 1380 3512
rect 1403 3507 1405 3512
rect 1429 3507 1431 3512
rect 425 3429 427 3434
rect 434 3429 436 3434
rect 239 3423 241 3428
rect 248 3423 250 3428
rect 281 3423 283 3428
rect 467 3429 469 3434
rect 555 3428 557 3433
rect 988 3436 990 3441
rect 997 3436 999 3441
rect 565 3428 567 3433
rect 611 3428 613 3433
rect 802 3430 804 3435
rect 811 3430 813 3435
rect 844 3430 846 3435
rect 1030 3436 1032 3441
rect 1118 3435 1120 3440
rect 1529 3508 1531 3513
rect 1555 3508 1557 3513
rect 1580 3508 1582 3513
rect 1606 3508 1608 3513
rect 1973 3538 1975 3543
rect 1999 3538 2001 3543
rect 2024 3538 2026 3543
rect 2050 3538 2052 3543
rect 2150 3539 2152 3544
rect 2176 3539 2178 3544
rect 2201 3539 2203 3544
rect 2227 3539 2229 3544
rect 1128 3435 1130 3440
rect 1174 3435 1176 3440
rect 1564 3422 1566 3427
rect 1573 3422 1575 3427
rect 1378 3416 1380 3421
rect 1387 3416 1389 3421
rect 1420 3416 1422 3421
rect 1606 3422 1608 3427
rect 1694 3421 1696 3426
rect 2185 3453 2187 3458
rect 2194 3453 2196 3458
rect 1999 3447 2001 3452
rect 2008 3447 2010 3452
rect 2041 3447 2043 3452
rect 2227 3453 2229 3458
rect 1704 3421 1706 3426
rect 1750 3421 1752 3426
rect 2315 3452 2317 3457
rect 2325 3452 2327 3457
rect 2371 3452 2373 3457
rect 400 3023 402 3028
rect 409 3023 411 3028
rect 442 3023 444 3028
rect 543 3023 545 3028
rect 552 3023 554 3028
rect 585 3023 587 3028
rect 706 3023 708 3028
rect 715 3023 717 3028
rect 748 3023 750 3028
rect 862 3023 864 3028
rect 871 3023 873 3028
rect 904 3023 906 3028
rect 1000 3023 1002 3028
rect 1009 3023 1011 3028
rect 1042 3023 1044 3028
rect 1143 3023 1145 3028
rect 1152 3023 1154 3028
rect 1185 3023 1187 3028
rect 1306 3023 1308 3028
rect 1315 3023 1317 3028
rect 1348 3023 1350 3028
rect 1462 3023 1464 3028
rect 1471 3023 1473 3028
rect 1504 3023 1506 3028
rect 2970 3214 2972 3219
rect 2996 3214 2998 3219
rect 3021 3214 3023 3219
rect 3047 3214 3049 3219
rect 3147 3215 3149 3220
rect 3173 3215 3175 3220
rect 3198 3215 3200 3220
rect 3224 3215 3226 3220
rect 3533 3221 3535 3226
rect 3559 3221 3561 3226
rect 3584 3221 3586 3226
rect 3610 3221 3612 3226
rect 3710 3222 3712 3227
rect 3736 3222 3738 3227
rect 3761 3222 3763 3227
rect 3787 3222 3789 3227
rect 4109 3207 4111 3212
rect 4135 3207 4137 3212
rect 4160 3207 4162 3212
rect 4186 3207 4188 3212
rect 3182 3129 3184 3134
rect 3191 3129 3193 3134
rect 2996 3123 2998 3128
rect 3005 3123 3007 3128
rect 3038 3123 3040 3128
rect 3224 3129 3226 3134
rect 3312 3128 3314 3133
rect 3745 3136 3747 3141
rect 3754 3136 3756 3141
rect 3322 3128 3324 3133
rect 3368 3128 3370 3133
rect 3559 3130 3561 3135
rect 3568 3130 3570 3135
rect 3601 3130 3603 3135
rect 3787 3136 3789 3141
rect 3875 3135 3877 3140
rect 4286 3208 4288 3213
rect 4312 3208 4314 3213
rect 4337 3208 4339 3213
rect 4363 3208 4365 3213
rect 4730 3238 4732 3243
rect 4756 3238 4758 3243
rect 4781 3238 4783 3243
rect 4807 3238 4809 3243
rect 4907 3239 4909 3244
rect 4933 3239 4935 3244
rect 4958 3239 4960 3244
rect 4984 3239 4986 3244
rect 3885 3135 3887 3140
rect 3931 3135 3933 3140
rect 4321 3122 4323 3127
rect 4330 3122 4332 3127
rect 4135 3116 4137 3121
rect 4144 3116 4146 3121
rect 4177 3116 4179 3121
rect 4363 3122 4365 3127
rect 4451 3121 4453 3126
rect 4942 3153 4944 3158
rect 4951 3153 4953 3158
rect 4756 3147 4758 3152
rect 4765 3147 4767 3152
rect 4798 3147 4800 3152
rect 4984 3153 4986 3158
rect 4461 3121 4463 3126
rect 4507 3121 4509 3126
rect 5072 3152 5074 3157
rect 5082 3152 5084 3157
rect 5128 3152 5130 3157
rect 242 2955 244 2960
rect 251 2955 253 2960
rect 284 2955 286 2960
rect 105 2871 107 2876
rect 114 2871 116 2876
rect 147 2871 149 2876
rect 194 2911 196 2915
rect 241 2874 243 2879
rect 250 2874 252 2879
rect 283 2874 285 2879
rect 400 2881 402 2886
rect 409 2881 411 2886
rect 442 2881 444 2886
rect 543 2881 545 2886
rect 552 2881 554 2886
rect 585 2881 587 2886
rect 706 2881 708 2886
rect 715 2881 717 2886
rect 748 2881 750 2886
rect 862 2881 864 2886
rect 871 2881 873 2886
rect 904 2881 906 2886
rect 1000 2881 1002 2886
rect 1009 2881 1011 2886
rect 1042 2881 1044 2886
rect 1143 2881 1145 2886
rect 1152 2881 1154 2886
rect 1185 2881 1187 2886
rect 1306 2881 1308 2886
rect 1315 2881 1317 2886
rect 1348 2881 1350 2886
rect 1462 2881 1464 2886
rect 1471 2881 1473 2886
rect 1504 2881 1506 2886
rect 1697 2904 1699 2909
rect 1723 2904 1725 2909
rect 1748 2904 1750 2909
rect 1774 2904 1776 2909
rect 1892 2905 1894 2910
rect 1918 2905 1920 2910
rect 1943 2905 1945 2910
rect 1969 2905 1971 2910
rect 2105 2904 2107 2909
rect 2131 2904 2133 2909
rect 2156 2904 2158 2909
rect 2182 2904 2184 2909
rect 2306 2905 2308 2910
rect 2332 2905 2334 2910
rect 2357 2905 2359 2910
rect 2383 2905 2385 2910
rect 194 2829 196 2833
rect 245 2783 247 2788
rect 254 2783 256 2788
rect 287 2783 289 2788
rect 400 2732 402 2737
rect 409 2732 411 2737
rect 442 2732 444 2737
rect 543 2732 545 2737
rect 552 2732 554 2737
rect 585 2732 587 2737
rect 706 2732 708 2737
rect 715 2732 717 2737
rect 748 2732 750 2737
rect 862 2732 864 2737
rect 871 2732 873 2737
rect 904 2732 906 2737
rect 1000 2732 1002 2737
rect 1009 2732 1011 2737
rect 1042 2732 1044 2737
rect 1143 2732 1145 2737
rect 1152 2732 1154 2737
rect 1185 2732 1187 2737
rect 1306 2732 1308 2737
rect 1315 2732 1317 2737
rect 1348 2732 1350 2737
rect 1462 2732 1464 2737
rect 1471 2732 1473 2737
rect 1504 2732 1506 2737
rect 2369 2707 2371 2717
rect 2384 2707 2386 2717
rect 2399 2707 2401 2717
rect 2414 2707 2416 2717
rect 2428 2707 2430 2717
rect 2454 2707 2456 2717
rect 400 2607 402 2612
rect 409 2607 411 2612
rect 442 2607 444 2612
rect 543 2607 545 2612
rect 552 2607 554 2612
rect 585 2607 587 2612
rect 706 2607 708 2612
rect 715 2607 717 2612
rect 748 2607 750 2612
rect 862 2607 864 2612
rect 871 2607 873 2612
rect 904 2607 906 2612
rect 1000 2607 1002 2612
rect 1009 2607 1011 2612
rect 1042 2607 1044 2612
rect 1143 2607 1145 2612
rect 1152 2607 1154 2612
rect 1185 2607 1187 2612
rect 1306 2607 1308 2612
rect 1315 2607 1317 2612
rect 1348 2607 1350 2612
rect 1462 2607 1464 2612
rect 1471 2607 1473 2612
rect 1504 2607 1506 2612
rect 782 2248 784 2253
rect 791 2248 793 2253
rect 824 2248 826 2253
rect 925 2248 927 2253
rect 934 2248 936 2253
rect 967 2248 969 2253
rect 1088 2248 1090 2253
rect 1097 2248 1099 2253
rect 1130 2248 1132 2253
rect 1244 2248 1246 2253
rect 1253 2248 1255 2253
rect 1286 2248 1288 2253
rect 2123 2664 2125 2668
rect 2818 2662 2820 2669
rect 2830 2662 2832 2669
rect 2845 2662 2847 2669
rect 2855 2662 2857 2669
rect 2878 2662 2880 2669
rect 2500 2607 2502 2617
rect 2515 2607 2517 2617
rect 2535 2607 2537 2617
rect 2545 2607 2547 2617
rect 2571 2607 2573 2617
rect 2125 2598 2127 2602
rect 2128 2531 2130 2535
rect 2128 2464 2130 2468
rect 2146 2359 2148 2363
rect 2046 2315 2048 2320
rect 2065 2315 2067 2320
rect 2090 2315 2092 2320
rect 2109 2315 2111 2320
rect 2148 2198 2150 2202
rect 2048 2154 2050 2159
rect 2067 2154 2069 2159
rect 2092 2154 2094 2159
rect 2111 2154 2113 2159
rect 2638 2569 2640 2579
rect 2653 2569 2655 2579
rect 2673 2569 2675 2579
rect 2697 2569 2699 2579
rect 2811 2541 2813 2545
rect 2764 2534 2766 2541
rect 2785 2534 2787 2541
rect 2747 2133 2749 2143
rect 2762 2133 2764 2143
rect 2782 2133 2784 2143
rect 2792 2133 2794 2143
rect 2818 2133 2820 2143
rect 2906 2133 2908 2138
rect 2917 2133 2919 2138
rect 2948 2133 2950 2138
rect 2147 2044 2149 2048
rect 2047 2000 2049 2005
rect 2066 2000 2068 2005
rect 2091 2000 2093 2005
rect 2110 2000 2112 2005
rect 2147 1896 2149 1900
rect 2809 1882 2811 1889
rect 2821 1882 2823 1889
rect 2836 1882 2838 1889
rect 2846 1882 2848 1889
rect 2869 1882 2871 1889
rect 2047 1852 2049 1857
rect 2066 1852 2068 1857
rect 2091 1852 2093 1857
rect 2110 1852 2112 1857
rect 2584 1818 2586 1828
rect 2599 1818 2601 1828
rect 2614 1818 2616 1828
rect 2629 1818 2631 1828
rect 2643 1818 2645 1828
rect 2669 1818 2671 1828
rect 2123 1769 2125 1773
rect 2452 1734 2454 1744
rect 2467 1734 2469 1744
rect 2487 1734 2489 1744
rect 2497 1734 2499 1744
rect 2523 1734 2525 1744
rect 2125 1703 2127 1707
rect 2311 1659 2313 1669
rect 2326 1659 2328 1669
rect 2346 1659 2348 1669
rect 2370 1659 2372 1669
rect 2128 1636 2130 1640
rect 2260 1597 2262 1601
rect 2213 1590 2215 1597
rect 2234 1590 2236 1597
rect 2128 1569 2130 1573
<< ptransistor >>
rect 213 3545 215 3550
rect 239 3545 241 3550
rect 264 3545 266 3550
rect 290 3545 292 3550
rect 390 3546 392 3551
rect 416 3546 418 3551
rect 441 3546 443 3551
rect 467 3546 469 3551
rect 776 3552 778 3557
rect 802 3552 804 3557
rect 827 3552 829 3557
rect 853 3552 855 3557
rect 239 3454 241 3459
rect 248 3454 250 3459
rect 281 3454 283 3459
rect 953 3553 955 3558
rect 979 3553 981 3558
rect 1004 3553 1006 3558
rect 1030 3553 1032 3558
rect 1352 3538 1354 3543
rect 1378 3538 1380 3543
rect 1403 3538 1405 3543
rect 1429 3538 1431 3543
rect 425 3460 427 3465
rect 434 3460 436 3465
rect 555 3467 557 3472
rect 565 3467 567 3472
rect 467 3460 469 3465
rect 611 3467 613 3472
rect 802 3461 804 3466
rect 811 3461 813 3466
rect 844 3461 846 3466
rect 988 3467 990 3472
rect 997 3467 999 3472
rect 1118 3474 1120 3479
rect 1128 3474 1130 3479
rect 1030 3467 1032 3472
rect 1174 3474 1176 3479
rect 1529 3539 1531 3544
rect 1555 3539 1557 3544
rect 1580 3539 1582 3544
rect 1606 3539 1608 3544
rect 1973 3569 1975 3574
rect 1999 3569 2001 3574
rect 2024 3569 2026 3574
rect 2050 3569 2052 3574
rect 2150 3570 2152 3575
rect 2176 3570 2178 3575
rect 2201 3570 2203 3575
rect 2227 3570 2229 3575
rect 1378 3447 1380 3452
rect 1387 3447 1389 3452
rect 1420 3447 1422 3452
rect 1564 3453 1566 3458
rect 1573 3453 1575 3458
rect 1694 3460 1696 3465
rect 1704 3460 1706 3465
rect 1606 3453 1608 3458
rect 1999 3478 2001 3483
rect 2008 3478 2010 3483
rect 2041 3478 2043 3483
rect 1750 3460 1752 3465
rect 2185 3484 2187 3489
rect 2194 3484 2196 3489
rect 2315 3491 2317 3496
rect 2325 3491 2327 3496
rect 2227 3484 2229 3489
rect 2371 3491 2373 3496
rect 400 3054 402 3059
rect 409 3054 411 3059
rect 442 3054 444 3059
rect 543 3054 545 3059
rect 552 3054 554 3059
rect 585 3054 587 3059
rect 706 3054 708 3059
rect 715 3054 717 3059
rect 748 3054 750 3059
rect 862 3054 864 3059
rect 871 3054 873 3059
rect 904 3054 906 3059
rect 1000 3054 1002 3059
rect 1009 3054 1011 3059
rect 1042 3054 1044 3059
rect 1143 3054 1145 3059
rect 1152 3054 1154 3059
rect 1185 3054 1187 3059
rect 1306 3054 1308 3059
rect 1315 3054 1317 3059
rect 1348 3054 1350 3059
rect 1462 3054 1464 3059
rect 1471 3054 1473 3059
rect 1504 3054 1506 3059
rect 2970 3245 2972 3250
rect 2996 3245 2998 3250
rect 3021 3245 3023 3250
rect 3047 3245 3049 3250
rect 3147 3246 3149 3251
rect 3173 3246 3175 3251
rect 3198 3246 3200 3251
rect 3224 3246 3226 3251
rect 3533 3252 3535 3257
rect 3559 3252 3561 3257
rect 3584 3252 3586 3257
rect 3610 3252 3612 3257
rect 2996 3154 2998 3159
rect 3005 3154 3007 3159
rect 3038 3154 3040 3159
rect 3710 3253 3712 3258
rect 3736 3253 3738 3258
rect 3761 3253 3763 3258
rect 3787 3253 3789 3258
rect 4109 3238 4111 3243
rect 4135 3238 4137 3243
rect 4160 3238 4162 3243
rect 4186 3238 4188 3243
rect 3182 3160 3184 3165
rect 3191 3160 3193 3165
rect 3312 3167 3314 3172
rect 3322 3167 3324 3172
rect 3224 3160 3226 3165
rect 3368 3167 3370 3172
rect 3559 3161 3561 3166
rect 3568 3161 3570 3166
rect 3601 3161 3603 3166
rect 3745 3167 3747 3172
rect 3754 3167 3756 3172
rect 3875 3174 3877 3179
rect 3885 3174 3887 3179
rect 3787 3167 3789 3172
rect 3931 3174 3933 3179
rect 4286 3239 4288 3244
rect 4312 3239 4314 3244
rect 4337 3239 4339 3244
rect 4363 3239 4365 3244
rect 4730 3269 4732 3274
rect 4756 3269 4758 3274
rect 4781 3269 4783 3274
rect 4807 3269 4809 3274
rect 4907 3270 4909 3275
rect 4933 3270 4935 3275
rect 4958 3270 4960 3275
rect 4984 3270 4986 3275
rect 4135 3147 4137 3152
rect 4144 3147 4146 3152
rect 4177 3147 4179 3152
rect 4321 3153 4323 3158
rect 4330 3153 4332 3158
rect 4451 3160 4453 3165
rect 4461 3160 4463 3165
rect 4363 3153 4365 3158
rect 4756 3178 4758 3183
rect 4765 3178 4767 3183
rect 4798 3178 4800 3183
rect 4507 3160 4509 3165
rect 4942 3184 4944 3189
rect 4951 3184 4953 3189
rect 5072 3191 5074 3196
rect 5082 3191 5084 3196
rect 4984 3184 4986 3189
rect 5128 3191 5130 3196
rect 242 2986 244 2991
rect 251 2986 253 2991
rect 284 2986 286 2991
rect 194 2934 196 2938
rect 105 2902 107 2907
rect 114 2902 116 2907
rect 147 2902 149 2907
rect 241 2905 243 2910
rect 250 2905 252 2910
rect 283 2905 285 2910
rect 194 2851 196 2855
rect 400 2912 402 2917
rect 409 2912 411 2917
rect 442 2912 444 2917
rect 543 2912 545 2917
rect 552 2912 554 2917
rect 585 2912 587 2917
rect 706 2912 708 2917
rect 715 2912 717 2917
rect 748 2912 750 2917
rect 862 2912 864 2917
rect 871 2912 873 2917
rect 904 2912 906 2917
rect 1000 2912 1002 2917
rect 1009 2912 1011 2917
rect 1042 2912 1044 2917
rect 1143 2912 1145 2917
rect 1152 2912 1154 2917
rect 1185 2912 1187 2917
rect 1306 2912 1308 2917
rect 1315 2912 1317 2917
rect 1348 2912 1350 2917
rect 1462 2912 1464 2917
rect 1471 2912 1473 2917
rect 1504 2912 1506 2917
rect 1697 2935 1699 2940
rect 1723 2935 1725 2940
rect 1748 2935 1750 2940
rect 1774 2935 1776 2940
rect 1892 2936 1894 2941
rect 1918 2936 1920 2941
rect 1943 2936 1945 2941
rect 1969 2936 1971 2941
rect 2105 2935 2107 2940
rect 2131 2935 2133 2940
rect 2156 2935 2158 2940
rect 2182 2935 2184 2940
rect 2306 2936 2308 2941
rect 2332 2936 2334 2941
rect 2357 2936 2359 2941
rect 2383 2936 2385 2941
rect 245 2814 247 2819
rect 254 2814 256 2819
rect 287 2814 289 2819
rect 400 2763 402 2768
rect 409 2763 411 2768
rect 442 2763 444 2768
rect 543 2763 545 2768
rect 552 2763 554 2768
rect 585 2763 587 2768
rect 706 2763 708 2768
rect 715 2763 717 2768
rect 748 2763 750 2768
rect 862 2763 864 2768
rect 871 2763 873 2768
rect 904 2763 906 2768
rect 1000 2763 1002 2768
rect 1009 2763 1011 2768
rect 1042 2763 1044 2768
rect 1143 2763 1145 2768
rect 1152 2763 1154 2768
rect 1185 2763 1187 2768
rect 1306 2763 1308 2768
rect 1315 2763 1317 2768
rect 1348 2763 1350 2768
rect 1462 2763 1464 2768
rect 1471 2763 1473 2768
rect 1504 2763 1506 2768
rect 2369 2742 2371 2752
rect 2384 2742 2386 2752
rect 2399 2742 2401 2752
rect 2414 2742 2416 2752
rect 2428 2742 2430 2752
rect 2454 2742 2456 2752
rect 2123 2688 2125 2692
rect 400 2638 402 2643
rect 409 2638 411 2643
rect 442 2638 444 2643
rect 543 2638 545 2643
rect 552 2638 554 2643
rect 585 2638 587 2643
rect 706 2638 708 2643
rect 715 2638 717 2643
rect 748 2638 750 2643
rect 862 2638 864 2643
rect 871 2638 873 2643
rect 904 2638 906 2643
rect 1000 2638 1002 2643
rect 1009 2638 1011 2643
rect 1042 2638 1044 2643
rect 1143 2638 1145 2643
rect 1152 2638 1154 2643
rect 1185 2638 1187 2643
rect 1306 2638 1308 2643
rect 1315 2638 1317 2643
rect 1348 2638 1350 2643
rect 1462 2638 1464 2643
rect 1471 2638 1473 2643
rect 1504 2638 1506 2643
rect 782 2279 784 2284
rect 791 2279 793 2284
rect 824 2279 826 2284
rect 925 2279 927 2284
rect 934 2279 936 2284
rect 967 2279 969 2284
rect 1088 2279 1090 2284
rect 1097 2279 1099 2284
rect 1130 2279 1132 2284
rect 1244 2279 1246 2284
rect 1253 2279 1255 2284
rect 1286 2279 1288 2284
rect 2500 2642 2502 2652
rect 2515 2642 2517 2652
rect 2535 2642 2537 2652
rect 2545 2642 2547 2652
rect 2571 2642 2573 2652
rect 2818 2692 2820 2699
rect 2830 2692 2832 2699
rect 2845 2692 2847 2699
rect 2855 2692 2857 2699
rect 2878 2692 2880 2699
rect 2125 2622 2127 2626
rect 2128 2555 2130 2559
rect 2128 2488 2130 2492
rect 2146 2383 2148 2387
rect 2046 2346 2048 2351
rect 2065 2346 2067 2351
rect 2090 2346 2092 2351
rect 2109 2346 2111 2351
rect 2148 2222 2150 2226
rect 2048 2185 2050 2190
rect 2067 2185 2069 2190
rect 2092 2185 2094 2190
rect 2111 2185 2113 2190
rect 2638 2604 2640 2614
rect 2653 2604 2655 2614
rect 2673 2604 2675 2614
rect 2697 2604 2699 2614
rect 2764 2564 2766 2569
rect 2785 2564 2787 2569
rect 2811 2565 2813 2569
rect 2747 2168 2749 2178
rect 2762 2168 2764 2178
rect 2782 2168 2784 2178
rect 2792 2168 2794 2178
rect 2818 2168 2820 2178
rect 2906 2164 2908 2169
rect 2917 2164 2919 2169
rect 2948 2164 2950 2169
rect 2147 2068 2149 2072
rect 2047 2031 2049 2036
rect 2066 2031 2068 2036
rect 2091 2031 2093 2036
rect 2110 2031 2112 2036
rect 2147 1920 2149 1924
rect 2809 1912 2811 1919
rect 2821 1912 2823 1919
rect 2836 1912 2838 1919
rect 2846 1912 2848 1919
rect 2869 1912 2871 1919
rect 2047 1883 2049 1888
rect 2066 1883 2068 1888
rect 2091 1883 2093 1888
rect 2110 1883 2112 1888
rect 2584 1853 2586 1863
rect 2599 1853 2601 1863
rect 2614 1853 2616 1863
rect 2629 1853 2631 1863
rect 2643 1853 2645 1863
rect 2669 1853 2671 1863
rect 2123 1793 2125 1797
rect 2452 1769 2454 1779
rect 2467 1769 2469 1779
rect 2487 1769 2489 1779
rect 2497 1769 2499 1779
rect 2523 1769 2525 1779
rect 2125 1727 2127 1731
rect 2311 1694 2313 1704
rect 2326 1694 2328 1704
rect 2346 1694 2348 1704
rect 2370 1694 2372 1704
rect 2128 1660 2130 1664
rect 2213 1620 2215 1625
rect 2234 1620 2236 1625
rect 2260 1621 2262 1625
rect 2128 1593 2130 1597
<< ndiffusion >>
rect 212 3515 213 3519
rect 208 3514 213 3515
rect 215 3515 217 3519
rect 215 3514 221 3515
rect 238 3515 239 3519
rect 234 3514 239 3515
rect 241 3515 243 3519
rect 241 3514 247 3515
rect 259 3518 264 3519
rect 263 3514 264 3518
rect 266 3515 269 3519
rect 266 3514 273 3515
rect 284 3518 290 3519
rect 288 3514 290 3518
rect 292 3515 293 3519
rect 292 3514 297 3515
rect 389 3516 390 3520
rect 385 3515 390 3516
rect 392 3516 394 3520
rect 392 3515 398 3516
rect 415 3516 416 3520
rect 411 3515 416 3516
rect 418 3516 420 3520
rect 418 3515 424 3516
rect 436 3519 441 3520
rect 440 3515 441 3519
rect 443 3516 446 3520
rect 443 3515 450 3516
rect 461 3519 467 3520
rect 465 3515 467 3519
rect 469 3516 470 3520
rect 469 3515 474 3516
rect 775 3522 776 3526
rect 771 3521 776 3522
rect 778 3522 780 3526
rect 778 3521 784 3522
rect 801 3522 802 3526
rect 797 3521 802 3522
rect 804 3522 806 3526
rect 804 3521 810 3522
rect 822 3525 827 3526
rect 826 3521 827 3525
rect 829 3522 832 3526
rect 829 3521 836 3522
rect 847 3525 853 3526
rect 851 3521 853 3525
rect 855 3522 856 3526
rect 855 3521 860 3522
rect 952 3523 953 3527
rect 948 3522 953 3523
rect 955 3523 957 3527
rect 955 3522 961 3523
rect 978 3523 979 3527
rect 974 3522 979 3523
rect 981 3523 983 3527
rect 981 3522 987 3523
rect 999 3526 1004 3527
rect 1003 3522 1004 3526
rect 1006 3523 1009 3527
rect 1006 3522 1013 3523
rect 1024 3526 1030 3527
rect 1028 3522 1030 3526
rect 1032 3523 1033 3527
rect 1032 3522 1037 3523
rect 1351 3508 1352 3512
rect 1347 3507 1352 3508
rect 1354 3508 1356 3512
rect 1354 3507 1360 3508
rect 1377 3508 1378 3512
rect 1373 3507 1378 3508
rect 1380 3508 1382 3512
rect 1380 3507 1386 3508
rect 1398 3511 1403 3512
rect 1402 3507 1403 3511
rect 1405 3508 1408 3512
rect 1405 3507 1412 3508
rect 1423 3511 1429 3512
rect 1427 3507 1429 3511
rect 1431 3508 1432 3512
rect 1431 3507 1436 3508
rect 420 3433 425 3434
rect 424 3429 425 3433
rect 427 3429 434 3434
rect 436 3430 438 3434
rect 436 3429 442 3430
rect 462 3432 467 3434
rect 234 3427 239 3428
rect 238 3423 239 3427
rect 241 3423 248 3428
rect 250 3424 252 3428
rect 250 3423 256 3424
rect 276 3426 281 3428
rect 280 3423 281 3426
rect 283 3425 286 3428
rect 466 3429 467 3432
rect 469 3431 472 3434
rect 469 3429 476 3431
rect 283 3423 290 3425
rect 550 3432 555 3433
rect 554 3428 555 3432
rect 557 3430 560 3433
rect 983 3440 988 3441
rect 987 3436 988 3440
rect 990 3436 997 3441
rect 999 3437 1001 3441
rect 999 3436 1005 3437
rect 1025 3439 1030 3441
rect 797 3434 802 3435
rect 564 3430 565 3433
rect 557 3428 565 3430
rect 567 3429 573 3433
rect 577 3429 585 3433
rect 567 3428 585 3429
rect 606 3431 611 3433
rect 610 3428 611 3431
rect 613 3430 616 3433
rect 801 3430 802 3434
rect 804 3430 811 3435
rect 813 3431 815 3435
rect 813 3430 819 3431
rect 839 3433 844 3435
rect 613 3428 620 3430
rect 843 3430 844 3433
rect 846 3432 849 3435
rect 1029 3436 1030 3439
rect 1032 3438 1035 3441
rect 1032 3436 1039 3438
rect 846 3430 853 3432
rect 1113 3439 1118 3440
rect 1117 3435 1118 3439
rect 1120 3437 1123 3440
rect 1528 3509 1529 3513
rect 1524 3508 1529 3509
rect 1531 3509 1533 3513
rect 1531 3508 1537 3509
rect 1554 3509 1555 3513
rect 1550 3508 1555 3509
rect 1557 3509 1559 3513
rect 1557 3508 1563 3509
rect 1575 3512 1580 3513
rect 1579 3508 1580 3512
rect 1582 3509 1585 3513
rect 1582 3508 1589 3509
rect 1600 3512 1606 3513
rect 1604 3508 1606 3512
rect 1608 3509 1609 3513
rect 1608 3508 1613 3509
rect 1972 3539 1973 3543
rect 1968 3538 1973 3539
rect 1975 3539 1977 3543
rect 1975 3538 1981 3539
rect 1998 3539 1999 3543
rect 1994 3538 1999 3539
rect 2001 3539 2003 3543
rect 2001 3538 2007 3539
rect 2019 3542 2024 3543
rect 2023 3538 2024 3542
rect 2026 3539 2029 3543
rect 2026 3538 2033 3539
rect 2044 3542 2050 3543
rect 2048 3538 2050 3542
rect 2052 3539 2053 3543
rect 2052 3538 2057 3539
rect 2149 3540 2150 3544
rect 2145 3539 2150 3540
rect 2152 3540 2154 3544
rect 2152 3539 2158 3540
rect 2175 3540 2176 3544
rect 2171 3539 2176 3540
rect 2178 3540 2180 3544
rect 2178 3539 2184 3540
rect 2196 3543 2201 3544
rect 2200 3539 2201 3543
rect 2203 3540 2206 3544
rect 2203 3539 2210 3540
rect 2221 3543 2227 3544
rect 2225 3539 2227 3543
rect 2229 3540 2230 3544
rect 2229 3539 2234 3540
rect 1127 3437 1128 3440
rect 1120 3435 1128 3437
rect 1130 3436 1136 3440
rect 1140 3436 1148 3440
rect 1130 3435 1148 3436
rect 1169 3438 1174 3440
rect 1173 3435 1174 3438
rect 1176 3437 1179 3440
rect 1176 3435 1183 3437
rect 1559 3426 1564 3427
rect 1563 3422 1564 3426
rect 1566 3422 1573 3427
rect 1575 3423 1577 3427
rect 1575 3422 1581 3423
rect 1601 3425 1606 3427
rect 1373 3420 1378 3421
rect 1377 3416 1378 3420
rect 1380 3416 1387 3421
rect 1389 3417 1391 3421
rect 1389 3416 1395 3417
rect 1415 3419 1420 3421
rect 1419 3416 1420 3419
rect 1422 3418 1425 3421
rect 1605 3422 1606 3425
rect 1608 3424 1611 3427
rect 1608 3422 1615 3424
rect 1422 3416 1429 3418
rect 1689 3425 1694 3426
rect 1693 3421 1694 3425
rect 1696 3423 1699 3426
rect 2180 3457 2185 3458
rect 2184 3453 2185 3457
rect 2187 3453 2194 3458
rect 2196 3454 2198 3458
rect 2196 3453 2202 3454
rect 2222 3456 2227 3458
rect 1994 3451 1999 3452
rect 1998 3447 1999 3451
rect 2001 3447 2008 3452
rect 2010 3448 2012 3452
rect 2010 3447 2016 3448
rect 2036 3450 2041 3452
rect 2040 3447 2041 3450
rect 2043 3449 2046 3452
rect 2226 3453 2227 3456
rect 2229 3455 2232 3458
rect 2229 3453 2236 3455
rect 2043 3447 2050 3449
rect 1703 3423 1704 3426
rect 1696 3421 1704 3423
rect 1706 3422 1712 3426
rect 1716 3422 1724 3426
rect 1706 3421 1724 3422
rect 1745 3424 1750 3426
rect 1749 3421 1750 3424
rect 1752 3423 1755 3426
rect 2310 3456 2315 3457
rect 2314 3452 2315 3456
rect 2317 3454 2320 3457
rect 2324 3454 2325 3457
rect 2317 3452 2325 3454
rect 2327 3453 2333 3457
rect 2337 3453 2345 3457
rect 2327 3452 2345 3453
rect 2366 3455 2371 3457
rect 2370 3452 2371 3455
rect 2373 3454 2376 3457
rect 2373 3452 2380 3454
rect 1752 3421 1759 3423
rect 395 3027 400 3028
rect 399 3023 400 3027
rect 402 3023 409 3028
rect 411 3024 413 3028
rect 411 3023 417 3024
rect 437 3026 442 3028
rect 441 3023 442 3026
rect 444 3025 447 3028
rect 444 3023 451 3025
rect 538 3027 543 3028
rect 542 3023 543 3027
rect 545 3023 552 3028
rect 554 3024 556 3028
rect 554 3023 560 3024
rect 580 3026 585 3028
rect 584 3023 585 3026
rect 587 3025 590 3028
rect 587 3023 594 3025
rect 701 3027 706 3028
rect 705 3023 706 3027
rect 708 3023 715 3028
rect 717 3024 719 3028
rect 717 3023 723 3024
rect 743 3026 748 3028
rect 747 3023 748 3026
rect 750 3025 753 3028
rect 750 3023 757 3025
rect 857 3027 862 3028
rect 861 3023 862 3027
rect 864 3023 871 3028
rect 873 3024 875 3028
rect 873 3023 879 3024
rect 899 3026 904 3028
rect 903 3023 904 3026
rect 906 3025 909 3028
rect 906 3023 913 3025
rect 995 3027 1000 3028
rect 999 3023 1000 3027
rect 1002 3023 1009 3028
rect 1011 3024 1013 3028
rect 1011 3023 1017 3024
rect 1037 3026 1042 3028
rect 1041 3023 1042 3026
rect 1044 3025 1047 3028
rect 1044 3023 1051 3025
rect 1138 3027 1143 3028
rect 1142 3023 1143 3027
rect 1145 3023 1152 3028
rect 1154 3024 1156 3028
rect 1154 3023 1160 3024
rect 1180 3026 1185 3028
rect 1184 3023 1185 3026
rect 1187 3025 1190 3028
rect 1187 3023 1194 3025
rect 1301 3027 1306 3028
rect 1305 3023 1306 3027
rect 1308 3023 1315 3028
rect 1317 3024 1319 3028
rect 1317 3023 1323 3024
rect 1343 3026 1348 3028
rect 1347 3023 1348 3026
rect 1350 3025 1353 3028
rect 1350 3023 1357 3025
rect 1457 3027 1462 3028
rect 1461 3023 1462 3027
rect 1464 3023 1471 3028
rect 1473 3024 1475 3028
rect 1473 3023 1479 3024
rect 1499 3026 1504 3028
rect 1503 3023 1504 3026
rect 1506 3025 1509 3028
rect 1506 3023 1513 3025
rect 2969 3215 2970 3219
rect 2965 3214 2970 3215
rect 2972 3215 2974 3219
rect 2972 3214 2978 3215
rect 2995 3215 2996 3219
rect 2991 3214 2996 3215
rect 2998 3215 3000 3219
rect 2998 3214 3004 3215
rect 3016 3218 3021 3219
rect 3020 3214 3021 3218
rect 3023 3215 3026 3219
rect 3023 3214 3030 3215
rect 3041 3218 3047 3219
rect 3045 3214 3047 3218
rect 3049 3215 3050 3219
rect 3049 3214 3054 3215
rect 3146 3216 3147 3220
rect 3142 3215 3147 3216
rect 3149 3216 3151 3220
rect 3149 3215 3155 3216
rect 3172 3216 3173 3220
rect 3168 3215 3173 3216
rect 3175 3216 3177 3220
rect 3175 3215 3181 3216
rect 3193 3219 3198 3220
rect 3197 3215 3198 3219
rect 3200 3216 3203 3220
rect 3200 3215 3207 3216
rect 3218 3219 3224 3220
rect 3222 3215 3224 3219
rect 3226 3216 3227 3220
rect 3226 3215 3231 3216
rect 3532 3222 3533 3226
rect 3528 3221 3533 3222
rect 3535 3222 3537 3226
rect 3535 3221 3541 3222
rect 3558 3222 3559 3226
rect 3554 3221 3559 3222
rect 3561 3222 3563 3226
rect 3561 3221 3567 3222
rect 3579 3225 3584 3226
rect 3583 3221 3584 3225
rect 3586 3222 3589 3226
rect 3586 3221 3593 3222
rect 3604 3225 3610 3226
rect 3608 3221 3610 3225
rect 3612 3222 3613 3226
rect 3612 3221 3617 3222
rect 3709 3223 3710 3227
rect 3705 3222 3710 3223
rect 3712 3223 3714 3227
rect 3712 3222 3718 3223
rect 3735 3223 3736 3227
rect 3731 3222 3736 3223
rect 3738 3223 3740 3227
rect 3738 3222 3744 3223
rect 3756 3226 3761 3227
rect 3760 3222 3761 3226
rect 3763 3223 3766 3227
rect 3763 3222 3770 3223
rect 3781 3226 3787 3227
rect 3785 3222 3787 3226
rect 3789 3223 3790 3227
rect 3789 3222 3794 3223
rect 4108 3208 4109 3212
rect 4104 3207 4109 3208
rect 4111 3208 4113 3212
rect 4111 3207 4117 3208
rect 4134 3208 4135 3212
rect 4130 3207 4135 3208
rect 4137 3208 4139 3212
rect 4137 3207 4143 3208
rect 4155 3211 4160 3212
rect 4159 3207 4160 3211
rect 4162 3208 4165 3212
rect 4162 3207 4169 3208
rect 4180 3211 4186 3212
rect 4184 3207 4186 3211
rect 4188 3208 4189 3212
rect 4188 3207 4193 3208
rect 3177 3133 3182 3134
rect 3181 3129 3182 3133
rect 3184 3129 3191 3134
rect 3193 3130 3195 3134
rect 3193 3129 3199 3130
rect 3219 3132 3224 3134
rect 2991 3127 2996 3128
rect 2995 3123 2996 3127
rect 2998 3123 3005 3128
rect 3007 3124 3009 3128
rect 3007 3123 3013 3124
rect 3033 3126 3038 3128
rect 3037 3123 3038 3126
rect 3040 3125 3043 3128
rect 3223 3129 3224 3132
rect 3226 3131 3229 3134
rect 3226 3129 3233 3131
rect 3040 3123 3047 3125
rect 3307 3132 3312 3133
rect 3311 3128 3312 3132
rect 3314 3130 3317 3133
rect 3740 3140 3745 3141
rect 3744 3136 3745 3140
rect 3747 3136 3754 3141
rect 3756 3137 3758 3141
rect 3756 3136 3762 3137
rect 3782 3139 3787 3141
rect 3554 3134 3559 3135
rect 3321 3130 3322 3133
rect 3314 3128 3322 3130
rect 3324 3129 3330 3133
rect 3334 3129 3342 3133
rect 3324 3128 3342 3129
rect 3363 3131 3368 3133
rect 3367 3128 3368 3131
rect 3370 3130 3373 3133
rect 3558 3130 3559 3134
rect 3561 3130 3568 3135
rect 3570 3131 3572 3135
rect 3570 3130 3576 3131
rect 3596 3133 3601 3135
rect 3370 3128 3377 3130
rect 3600 3130 3601 3133
rect 3603 3132 3606 3135
rect 3786 3136 3787 3139
rect 3789 3138 3792 3141
rect 3789 3136 3796 3138
rect 3603 3130 3610 3132
rect 3870 3139 3875 3140
rect 3874 3135 3875 3139
rect 3877 3137 3880 3140
rect 4285 3209 4286 3213
rect 4281 3208 4286 3209
rect 4288 3209 4290 3213
rect 4288 3208 4294 3209
rect 4311 3209 4312 3213
rect 4307 3208 4312 3209
rect 4314 3209 4316 3213
rect 4314 3208 4320 3209
rect 4332 3212 4337 3213
rect 4336 3208 4337 3212
rect 4339 3209 4342 3213
rect 4339 3208 4346 3209
rect 4357 3212 4363 3213
rect 4361 3208 4363 3212
rect 4365 3209 4366 3213
rect 4365 3208 4370 3209
rect 4729 3239 4730 3243
rect 4725 3238 4730 3239
rect 4732 3239 4734 3243
rect 4732 3238 4738 3239
rect 4755 3239 4756 3243
rect 4751 3238 4756 3239
rect 4758 3239 4760 3243
rect 4758 3238 4764 3239
rect 4776 3242 4781 3243
rect 4780 3238 4781 3242
rect 4783 3239 4786 3243
rect 4783 3238 4790 3239
rect 4801 3242 4807 3243
rect 4805 3238 4807 3242
rect 4809 3239 4810 3243
rect 4809 3238 4814 3239
rect 4906 3240 4907 3244
rect 4902 3239 4907 3240
rect 4909 3240 4911 3244
rect 4909 3239 4915 3240
rect 4932 3240 4933 3244
rect 4928 3239 4933 3240
rect 4935 3240 4937 3244
rect 4935 3239 4941 3240
rect 4953 3243 4958 3244
rect 4957 3239 4958 3243
rect 4960 3240 4963 3244
rect 4960 3239 4967 3240
rect 4978 3243 4984 3244
rect 4982 3239 4984 3243
rect 4986 3240 4987 3244
rect 4986 3239 4991 3240
rect 3884 3137 3885 3140
rect 3877 3135 3885 3137
rect 3887 3136 3893 3140
rect 3897 3136 3905 3140
rect 3887 3135 3905 3136
rect 3926 3138 3931 3140
rect 3930 3135 3931 3138
rect 3933 3137 3936 3140
rect 3933 3135 3940 3137
rect 4316 3126 4321 3127
rect 4320 3122 4321 3126
rect 4323 3122 4330 3127
rect 4332 3123 4334 3127
rect 4332 3122 4338 3123
rect 4358 3125 4363 3127
rect 4130 3120 4135 3121
rect 4134 3116 4135 3120
rect 4137 3116 4144 3121
rect 4146 3117 4148 3121
rect 4146 3116 4152 3117
rect 4172 3119 4177 3121
rect 4176 3116 4177 3119
rect 4179 3118 4182 3121
rect 4362 3122 4363 3125
rect 4365 3124 4368 3127
rect 4365 3122 4372 3124
rect 4179 3116 4186 3118
rect 4446 3125 4451 3126
rect 4450 3121 4451 3125
rect 4453 3123 4456 3126
rect 4937 3157 4942 3158
rect 4941 3153 4942 3157
rect 4944 3153 4951 3158
rect 4953 3154 4955 3158
rect 4953 3153 4959 3154
rect 4979 3156 4984 3158
rect 4751 3151 4756 3152
rect 4755 3147 4756 3151
rect 4758 3147 4765 3152
rect 4767 3148 4769 3152
rect 4767 3147 4773 3148
rect 4793 3150 4798 3152
rect 4797 3147 4798 3150
rect 4800 3149 4803 3152
rect 4983 3153 4984 3156
rect 4986 3155 4989 3158
rect 4986 3153 4993 3155
rect 4800 3147 4807 3149
rect 4460 3123 4461 3126
rect 4453 3121 4461 3123
rect 4463 3122 4469 3126
rect 4473 3122 4481 3126
rect 4463 3121 4481 3122
rect 4502 3124 4507 3126
rect 4506 3121 4507 3124
rect 4509 3123 4512 3126
rect 5067 3156 5072 3157
rect 5071 3152 5072 3156
rect 5074 3154 5077 3157
rect 5081 3154 5082 3157
rect 5074 3152 5082 3154
rect 5084 3153 5090 3157
rect 5094 3153 5102 3157
rect 5084 3152 5102 3153
rect 5123 3155 5128 3157
rect 5127 3152 5128 3155
rect 5130 3154 5133 3157
rect 5130 3152 5137 3154
rect 4509 3121 4516 3123
rect 237 2959 242 2960
rect 241 2955 242 2959
rect 244 2955 251 2960
rect 253 2956 255 2960
rect 253 2955 259 2956
rect 279 2958 284 2960
rect 283 2955 284 2958
rect 286 2957 289 2960
rect 286 2955 293 2957
rect 100 2875 105 2876
rect 104 2871 105 2875
rect 107 2871 114 2876
rect 116 2872 118 2876
rect 116 2871 122 2872
rect 142 2874 147 2876
rect 146 2871 147 2874
rect 149 2873 152 2876
rect 149 2871 156 2873
rect 193 2911 194 2915
rect 196 2911 197 2915
rect 236 2878 241 2879
rect 240 2874 241 2878
rect 243 2874 250 2879
rect 252 2875 254 2879
rect 252 2874 258 2875
rect 278 2877 283 2879
rect 282 2874 283 2877
rect 285 2876 288 2879
rect 285 2874 292 2876
rect 395 2885 400 2886
rect 399 2881 400 2885
rect 402 2881 409 2886
rect 411 2882 413 2886
rect 411 2881 417 2882
rect 437 2884 442 2886
rect 441 2881 442 2884
rect 444 2883 447 2886
rect 444 2881 451 2883
rect 538 2885 543 2886
rect 542 2881 543 2885
rect 545 2881 552 2886
rect 554 2882 556 2886
rect 554 2881 560 2882
rect 580 2884 585 2886
rect 584 2881 585 2884
rect 587 2883 590 2886
rect 587 2881 594 2883
rect 701 2885 706 2886
rect 705 2881 706 2885
rect 708 2881 715 2886
rect 717 2882 719 2886
rect 717 2881 723 2882
rect 743 2884 748 2886
rect 747 2881 748 2884
rect 750 2883 753 2886
rect 750 2881 757 2883
rect 857 2885 862 2886
rect 861 2881 862 2885
rect 864 2881 871 2886
rect 873 2882 875 2886
rect 873 2881 879 2882
rect 899 2884 904 2886
rect 903 2881 904 2884
rect 906 2883 909 2886
rect 906 2881 913 2883
rect 995 2885 1000 2886
rect 999 2881 1000 2885
rect 1002 2881 1009 2886
rect 1011 2882 1013 2886
rect 1011 2881 1017 2882
rect 1037 2884 1042 2886
rect 1041 2881 1042 2884
rect 1044 2883 1047 2886
rect 1044 2881 1051 2883
rect 1138 2885 1143 2886
rect 1142 2881 1143 2885
rect 1145 2881 1152 2886
rect 1154 2882 1156 2886
rect 1154 2881 1160 2882
rect 1180 2884 1185 2886
rect 1184 2881 1185 2884
rect 1187 2883 1190 2886
rect 1187 2881 1194 2883
rect 1301 2885 1306 2886
rect 1305 2881 1306 2885
rect 1308 2881 1315 2886
rect 1317 2882 1319 2886
rect 1317 2881 1323 2882
rect 1343 2884 1348 2886
rect 1347 2881 1348 2884
rect 1350 2883 1353 2886
rect 1350 2881 1357 2883
rect 1457 2885 1462 2886
rect 1461 2881 1462 2885
rect 1464 2881 1471 2886
rect 1473 2882 1475 2886
rect 1473 2881 1479 2882
rect 1499 2884 1504 2886
rect 1503 2881 1504 2884
rect 1506 2883 1509 2886
rect 1506 2881 1513 2883
rect 1696 2905 1697 2909
rect 1692 2904 1697 2905
rect 1699 2905 1701 2909
rect 1699 2904 1705 2905
rect 1722 2905 1723 2909
rect 1718 2904 1723 2905
rect 1725 2905 1727 2909
rect 1725 2904 1731 2905
rect 1743 2908 1748 2909
rect 1747 2904 1748 2908
rect 1750 2905 1753 2909
rect 1750 2904 1757 2905
rect 1768 2908 1774 2909
rect 1772 2904 1774 2908
rect 1776 2905 1777 2909
rect 1776 2904 1781 2905
rect 1891 2906 1892 2910
rect 1887 2905 1892 2906
rect 1894 2906 1896 2910
rect 1894 2905 1900 2906
rect 1917 2906 1918 2910
rect 1913 2905 1918 2906
rect 1920 2906 1922 2910
rect 1920 2905 1926 2906
rect 1938 2909 1943 2910
rect 1942 2905 1943 2909
rect 1945 2906 1948 2910
rect 1945 2905 1952 2906
rect 1963 2909 1969 2910
rect 1967 2905 1969 2909
rect 1971 2906 1972 2910
rect 1971 2905 1976 2906
rect 2104 2905 2105 2909
rect 2100 2904 2105 2905
rect 2107 2905 2109 2909
rect 2107 2904 2113 2905
rect 2130 2905 2131 2909
rect 2126 2904 2131 2905
rect 2133 2905 2135 2909
rect 2133 2904 2139 2905
rect 2151 2908 2156 2909
rect 2155 2904 2156 2908
rect 2158 2905 2161 2909
rect 2158 2904 2165 2905
rect 2176 2908 2182 2909
rect 2180 2904 2182 2908
rect 2184 2905 2185 2909
rect 2184 2904 2189 2905
rect 2305 2906 2306 2910
rect 2301 2905 2306 2906
rect 2308 2906 2310 2910
rect 2308 2905 2314 2906
rect 2331 2906 2332 2910
rect 2327 2905 2332 2906
rect 2334 2906 2336 2910
rect 2334 2905 2340 2906
rect 2352 2909 2357 2910
rect 2356 2905 2357 2909
rect 2359 2906 2362 2910
rect 2359 2905 2366 2906
rect 2377 2909 2383 2910
rect 2381 2905 2383 2909
rect 2385 2906 2386 2910
rect 2385 2905 2390 2906
rect 193 2829 194 2833
rect 196 2829 197 2833
rect 240 2787 245 2788
rect 244 2783 245 2787
rect 247 2783 254 2788
rect 256 2784 258 2788
rect 256 2783 262 2784
rect 282 2786 287 2788
rect 286 2783 287 2786
rect 289 2785 292 2788
rect 289 2783 296 2785
rect 395 2736 400 2737
rect 399 2732 400 2736
rect 402 2732 409 2737
rect 411 2733 413 2737
rect 411 2732 417 2733
rect 437 2735 442 2737
rect 441 2732 442 2735
rect 444 2734 447 2737
rect 444 2732 451 2734
rect 538 2736 543 2737
rect 542 2732 543 2736
rect 545 2732 552 2737
rect 554 2733 556 2737
rect 554 2732 560 2733
rect 580 2735 585 2737
rect 584 2732 585 2735
rect 587 2734 590 2737
rect 587 2732 594 2734
rect 701 2736 706 2737
rect 705 2732 706 2736
rect 708 2732 715 2737
rect 717 2733 719 2737
rect 717 2732 723 2733
rect 743 2735 748 2737
rect 747 2732 748 2735
rect 750 2734 753 2737
rect 750 2732 757 2734
rect 857 2736 862 2737
rect 861 2732 862 2736
rect 864 2732 871 2737
rect 873 2733 875 2737
rect 873 2732 879 2733
rect 899 2735 904 2737
rect 903 2732 904 2735
rect 906 2734 909 2737
rect 906 2732 913 2734
rect 995 2736 1000 2737
rect 999 2732 1000 2736
rect 1002 2732 1009 2737
rect 1011 2733 1013 2737
rect 1011 2732 1017 2733
rect 1037 2735 1042 2737
rect 1041 2732 1042 2735
rect 1044 2734 1047 2737
rect 1044 2732 1051 2734
rect 1138 2736 1143 2737
rect 1142 2732 1143 2736
rect 1145 2732 1152 2737
rect 1154 2733 1156 2737
rect 1154 2732 1160 2733
rect 1180 2735 1185 2737
rect 1184 2732 1185 2735
rect 1187 2734 1190 2737
rect 1187 2732 1194 2734
rect 1301 2736 1306 2737
rect 1305 2732 1306 2736
rect 1308 2732 1315 2737
rect 1317 2733 1319 2737
rect 1317 2732 1323 2733
rect 1343 2735 1348 2737
rect 1347 2732 1348 2735
rect 1350 2734 1353 2737
rect 1350 2732 1357 2734
rect 1457 2736 1462 2737
rect 1461 2732 1462 2736
rect 1464 2732 1471 2737
rect 1473 2733 1475 2737
rect 1473 2732 1479 2733
rect 1499 2735 1504 2737
rect 1503 2732 1504 2735
rect 1506 2734 1509 2737
rect 1506 2732 1513 2734
rect 2360 2711 2369 2717
rect 2364 2707 2369 2711
rect 2371 2707 2384 2717
rect 2386 2707 2399 2717
rect 2401 2707 2414 2717
rect 2416 2707 2428 2717
rect 2430 2711 2439 2717
rect 2430 2707 2435 2711
rect 2445 2711 2454 2717
rect 2449 2707 2454 2711
rect 2456 2713 2461 2717
rect 2456 2707 2465 2713
rect 395 2611 400 2612
rect 399 2607 400 2611
rect 402 2607 409 2612
rect 411 2608 413 2612
rect 411 2607 417 2608
rect 437 2610 442 2612
rect 441 2607 442 2610
rect 444 2609 447 2612
rect 444 2607 451 2609
rect 538 2611 543 2612
rect 542 2607 543 2611
rect 545 2607 552 2612
rect 554 2608 556 2612
rect 554 2607 560 2608
rect 580 2610 585 2612
rect 584 2607 585 2610
rect 587 2609 590 2612
rect 587 2607 594 2609
rect 701 2611 706 2612
rect 705 2607 706 2611
rect 708 2607 715 2612
rect 717 2608 719 2612
rect 717 2607 723 2608
rect 743 2610 748 2612
rect 747 2607 748 2610
rect 750 2609 753 2612
rect 750 2607 757 2609
rect 857 2611 862 2612
rect 861 2607 862 2611
rect 864 2607 871 2612
rect 873 2608 875 2612
rect 873 2607 879 2608
rect 899 2610 904 2612
rect 903 2607 904 2610
rect 906 2609 909 2612
rect 906 2607 913 2609
rect 995 2611 1000 2612
rect 999 2607 1000 2611
rect 1002 2607 1009 2612
rect 1011 2608 1013 2612
rect 1011 2607 1017 2608
rect 1037 2610 1042 2612
rect 1041 2607 1042 2610
rect 1044 2609 1047 2612
rect 1044 2607 1051 2609
rect 1138 2611 1143 2612
rect 1142 2607 1143 2611
rect 1145 2607 1152 2612
rect 1154 2608 1156 2612
rect 1154 2607 1160 2608
rect 1180 2610 1185 2612
rect 1184 2607 1185 2610
rect 1187 2609 1190 2612
rect 1187 2607 1194 2609
rect 1301 2611 1306 2612
rect 1305 2607 1306 2611
rect 1308 2607 1315 2612
rect 1317 2608 1319 2612
rect 1317 2607 1323 2608
rect 1343 2610 1348 2612
rect 1347 2607 1348 2610
rect 1350 2609 1353 2612
rect 1350 2607 1357 2609
rect 1457 2611 1462 2612
rect 1461 2607 1462 2611
rect 1464 2607 1471 2612
rect 1473 2608 1475 2612
rect 1473 2607 1479 2608
rect 1499 2610 1504 2612
rect 1503 2607 1504 2610
rect 1506 2609 1509 2612
rect 1506 2607 1513 2609
rect 777 2252 782 2253
rect 781 2248 782 2252
rect 784 2248 791 2253
rect 793 2249 795 2253
rect 793 2248 799 2249
rect 819 2251 824 2253
rect 823 2248 824 2251
rect 826 2250 829 2253
rect 826 2248 833 2250
rect 920 2252 925 2253
rect 924 2248 925 2252
rect 927 2248 934 2253
rect 936 2249 938 2253
rect 936 2248 942 2249
rect 962 2251 967 2253
rect 966 2248 967 2251
rect 969 2250 972 2253
rect 969 2248 976 2250
rect 1083 2252 1088 2253
rect 1087 2248 1088 2252
rect 1090 2248 1097 2253
rect 1099 2249 1101 2253
rect 1099 2248 1105 2249
rect 1125 2251 1130 2253
rect 1129 2248 1130 2251
rect 1132 2250 1135 2253
rect 1132 2248 1139 2250
rect 1239 2252 1244 2253
rect 1243 2248 1244 2252
rect 1246 2248 1253 2253
rect 1255 2249 1257 2253
rect 1255 2248 1261 2249
rect 1281 2251 1286 2253
rect 1285 2248 1286 2251
rect 1288 2250 1291 2253
rect 1288 2248 1295 2250
rect 2122 2664 2123 2668
rect 2125 2664 2126 2668
rect 2810 2666 2818 2669
rect 2814 2662 2818 2666
rect 2820 2665 2823 2669
rect 2827 2665 2830 2669
rect 2820 2662 2830 2665
rect 2832 2666 2845 2669
rect 2832 2662 2836 2666
rect 2840 2662 2845 2666
rect 2847 2665 2849 2669
rect 2853 2665 2855 2669
rect 2847 2662 2855 2665
rect 2857 2665 2862 2669
rect 2857 2662 2866 2665
rect 2874 2665 2878 2669
rect 2870 2662 2878 2665
rect 2880 2665 2883 2669
rect 2880 2662 2887 2665
rect 2491 2611 2500 2617
rect 2495 2607 2500 2611
rect 2502 2607 2515 2617
rect 2517 2607 2535 2617
rect 2537 2607 2545 2617
rect 2547 2611 2557 2617
rect 2547 2607 2553 2611
rect 2562 2611 2571 2617
rect 2566 2607 2571 2611
rect 2573 2613 2578 2617
rect 2573 2607 2582 2613
rect 2124 2598 2125 2602
rect 2127 2598 2128 2602
rect 2127 2531 2128 2535
rect 2130 2531 2131 2535
rect 2127 2464 2128 2468
rect 2130 2464 2131 2468
rect 2145 2359 2146 2363
rect 2148 2359 2149 2363
rect 2041 2319 2046 2320
rect 2045 2315 2046 2319
rect 2048 2319 2052 2320
rect 2060 2319 2065 2320
rect 2048 2315 2050 2319
rect 2064 2315 2065 2319
rect 2067 2319 2073 2320
rect 2067 2315 2069 2319
rect 2085 2319 2090 2320
rect 2089 2315 2090 2319
rect 2092 2319 2098 2320
rect 2092 2315 2094 2319
rect 2104 2319 2109 2320
rect 2108 2315 2109 2319
rect 2111 2319 2117 2320
rect 2111 2315 2113 2319
rect 2147 2198 2148 2202
rect 2150 2198 2151 2202
rect 2043 2158 2048 2159
rect 2047 2154 2048 2158
rect 2050 2158 2054 2159
rect 2062 2158 2067 2159
rect 2050 2154 2052 2158
rect 2066 2154 2067 2158
rect 2069 2158 2075 2159
rect 2069 2154 2071 2158
rect 2087 2158 2092 2159
rect 2091 2154 2092 2158
rect 2094 2158 2100 2159
rect 2094 2154 2096 2158
rect 2106 2158 2111 2159
rect 2110 2154 2111 2158
rect 2113 2158 2119 2159
rect 2113 2154 2115 2158
rect 2629 2573 2638 2579
rect 2633 2569 2638 2573
rect 2640 2569 2653 2579
rect 2655 2569 2673 2579
rect 2675 2573 2683 2579
rect 2675 2569 2679 2573
rect 2688 2573 2697 2579
rect 2692 2569 2697 2573
rect 2699 2575 2704 2579
rect 2699 2569 2708 2575
rect 2810 2541 2811 2545
rect 2813 2541 2814 2545
rect 2762 2537 2764 2541
rect 2758 2534 2764 2537
rect 2766 2534 2785 2541
rect 2787 2538 2794 2541
rect 2787 2534 2790 2538
rect 2738 2137 2747 2143
rect 2742 2133 2747 2137
rect 2749 2133 2762 2143
rect 2764 2133 2782 2143
rect 2784 2133 2792 2143
rect 2794 2137 2804 2143
rect 2794 2133 2800 2137
rect 2809 2137 2818 2143
rect 2813 2133 2818 2137
rect 2820 2139 2825 2143
rect 2820 2133 2829 2139
rect 2901 2137 2906 2138
rect 2905 2133 2906 2137
rect 2908 2133 2917 2138
rect 2919 2134 2920 2138
rect 2919 2133 2924 2134
rect 2943 2136 2948 2138
rect 2947 2133 2948 2136
rect 2950 2135 2953 2138
rect 2950 2133 2957 2135
rect 2146 2044 2147 2048
rect 2149 2044 2150 2048
rect 2042 2004 2047 2005
rect 2046 2000 2047 2004
rect 2049 2004 2053 2005
rect 2061 2004 2066 2005
rect 2049 2000 2051 2004
rect 2065 2000 2066 2004
rect 2068 2004 2074 2005
rect 2068 2000 2070 2004
rect 2086 2004 2091 2005
rect 2090 2000 2091 2004
rect 2093 2004 2099 2005
rect 2093 2000 2095 2004
rect 2105 2004 2110 2005
rect 2109 2000 2110 2004
rect 2112 2004 2118 2005
rect 2112 2000 2114 2004
rect 2146 1896 2147 1900
rect 2149 1896 2150 1900
rect 2801 1886 2809 1889
rect 2805 1882 2809 1886
rect 2811 1885 2814 1889
rect 2818 1885 2821 1889
rect 2811 1882 2821 1885
rect 2823 1886 2836 1889
rect 2823 1882 2827 1886
rect 2831 1882 2836 1886
rect 2838 1885 2840 1889
rect 2844 1885 2846 1889
rect 2838 1882 2846 1885
rect 2848 1885 2853 1889
rect 2848 1882 2857 1885
rect 2865 1885 2869 1889
rect 2861 1882 2869 1885
rect 2871 1885 2874 1889
rect 2871 1882 2878 1885
rect 2042 1856 2047 1857
rect 2046 1852 2047 1856
rect 2049 1856 2053 1857
rect 2061 1856 2066 1857
rect 2049 1852 2051 1856
rect 2065 1852 2066 1856
rect 2068 1856 2074 1857
rect 2068 1852 2070 1856
rect 2086 1856 2091 1857
rect 2090 1852 2091 1856
rect 2093 1856 2099 1857
rect 2093 1852 2095 1856
rect 2105 1856 2110 1857
rect 2109 1852 2110 1856
rect 2112 1856 2118 1857
rect 2112 1852 2114 1856
rect 2575 1822 2584 1828
rect 2579 1818 2584 1822
rect 2586 1818 2599 1828
rect 2601 1818 2614 1828
rect 2616 1818 2629 1828
rect 2631 1818 2643 1828
rect 2645 1822 2654 1828
rect 2645 1818 2650 1822
rect 2660 1822 2669 1828
rect 2664 1818 2669 1822
rect 2671 1824 2676 1828
rect 2671 1818 2680 1824
rect 2122 1769 2123 1773
rect 2125 1769 2126 1773
rect 2443 1738 2452 1744
rect 2447 1734 2452 1738
rect 2454 1734 2467 1744
rect 2469 1734 2487 1744
rect 2489 1734 2497 1744
rect 2499 1738 2509 1744
rect 2499 1734 2505 1738
rect 2514 1738 2523 1744
rect 2518 1734 2523 1738
rect 2525 1740 2530 1744
rect 2525 1734 2534 1740
rect 2124 1703 2125 1707
rect 2127 1703 2128 1707
rect 2302 1663 2311 1669
rect 2306 1659 2311 1663
rect 2313 1659 2326 1669
rect 2328 1659 2346 1669
rect 2348 1663 2356 1669
rect 2348 1659 2352 1663
rect 2361 1663 2370 1669
rect 2365 1659 2370 1663
rect 2372 1665 2377 1669
rect 2372 1659 2381 1665
rect 2127 1636 2128 1640
rect 2130 1636 2131 1640
rect 2259 1597 2260 1601
rect 2262 1597 2263 1601
rect 2211 1593 2213 1597
rect 2207 1590 2213 1593
rect 2215 1590 2234 1597
rect 2236 1594 2243 1597
rect 2236 1590 2239 1594
rect 2127 1569 2128 1573
rect 2130 1569 2131 1573
<< pdiffusion >>
rect 208 3549 213 3550
rect 212 3545 213 3549
rect 215 3549 221 3550
rect 215 3545 217 3549
rect 234 3549 239 3550
rect 238 3545 239 3549
rect 241 3549 247 3550
rect 241 3545 243 3549
rect 263 3546 264 3550
rect 259 3545 264 3546
rect 266 3549 273 3550
rect 266 3545 269 3549
rect 288 3547 290 3550
rect 284 3545 290 3547
rect 292 3549 297 3550
rect 292 3545 293 3549
rect 385 3550 390 3551
rect 389 3546 390 3550
rect 392 3550 398 3551
rect 392 3546 394 3550
rect 411 3550 416 3551
rect 415 3546 416 3550
rect 418 3550 424 3551
rect 418 3546 420 3550
rect 440 3547 441 3551
rect 436 3546 441 3547
rect 443 3550 450 3551
rect 443 3546 446 3550
rect 465 3548 467 3551
rect 461 3546 467 3548
rect 469 3550 474 3551
rect 469 3546 470 3550
rect 771 3556 776 3557
rect 775 3552 776 3556
rect 778 3556 784 3557
rect 778 3552 780 3556
rect 797 3556 802 3557
rect 801 3552 802 3556
rect 804 3556 810 3557
rect 804 3552 806 3556
rect 826 3553 827 3557
rect 822 3552 827 3553
rect 829 3556 836 3557
rect 829 3552 832 3556
rect 851 3554 853 3557
rect 847 3552 853 3554
rect 855 3556 860 3557
rect 855 3552 856 3556
rect 238 3456 239 3459
rect 234 3454 239 3456
rect 241 3457 248 3459
rect 241 3454 243 3457
rect 247 3454 248 3457
rect 250 3456 252 3459
rect 250 3454 256 3456
rect 280 3456 281 3459
rect 276 3454 281 3456
rect 283 3455 286 3459
rect 283 3454 290 3455
rect 948 3557 953 3558
rect 952 3553 953 3557
rect 955 3557 961 3558
rect 955 3553 957 3557
rect 974 3557 979 3558
rect 978 3553 979 3557
rect 981 3557 987 3558
rect 981 3553 983 3557
rect 1003 3554 1004 3558
rect 999 3553 1004 3554
rect 1006 3557 1013 3558
rect 1006 3553 1009 3557
rect 1028 3555 1030 3558
rect 1024 3553 1030 3555
rect 1032 3557 1037 3558
rect 1032 3553 1033 3557
rect 1347 3542 1352 3543
rect 1351 3538 1352 3542
rect 1354 3542 1360 3543
rect 1354 3538 1356 3542
rect 1373 3542 1378 3543
rect 1377 3538 1378 3542
rect 1380 3542 1386 3543
rect 1380 3538 1382 3542
rect 1402 3539 1403 3543
rect 1398 3538 1403 3539
rect 1405 3542 1412 3543
rect 1405 3538 1408 3542
rect 1427 3540 1429 3543
rect 1423 3538 1429 3540
rect 1431 3542 1436 3543
rect 1431 3538 1432 3542
rect 554 3469 555 3472
rect 424 3462 425 3465
rect 420 3460 425 3462
rect 427 3463 434 3465
rect 427 3460 429 3463
rect 433 3460 434 3463
rect 436 3462 438 3465
rect 436 3460 442 3462
rect 550 3467 555 3469
rect 557 3467 565 3472
rect 567 3470 585 3472
rect 567 3467 573 3470
rect 466 3462 467 3465
rect 462 3460 467 3462
rect 469 3461 472 3465
rect 469 3460 476 3461
rect 577 3467 585 3470
rect 610 3469 611 3472
rect 606 3467 611 3469
rect 613 3468 616 3472
rect 613 3467 620 3468
rect 801 3463 802 3466
rect 797 3461 802 3463
rect 804 3464 811 3466
rect 804 3461 806 3464
rect 810 3461 811 3464
rect 813 3463 815 3466
rect 813 3461 819 3463
rect 843 3463 844 3466
rect 839 3461 844 3463
rect 846 3462 849 3466
rect 846 3461 853 3462
rect 1117 3476 1118 3479
rect 987 3469 988 3472
rect 983 3467 988 3469
rect 990 3470 997 3472
rect 990 3467 992 3470
rect 996 3467 997 3470
rect 999 3469 1001 3472
rect 999 3467 1005 3469
rect 1113 3474 1118 3476
rect 1120 3474 1128 3479
rect 1130 3477 1148 3479
rect 1130 3474 1136 3477
rect 1029 3469 1030 3472
rect 1025 3467 1030 3469
rect 1032 3468 1035 3472
rect 1032 3467 1039 3468
rect 1140 3474 1148 3477
rect 1173 3476 1174 3479
rect 1169 3474 1174 3476
rect 1176 3475 1179 3479
rect 1176 3474 1183 3475
rect 1524 3543 1529 3544
rect 1528 3539 1529 3543
rect 1531 3543 1537 3544
rect 1531 3539 1533 3543
rect 1550 3543 1555 3544
rect 1554 3539 1555 3543
rect 1557 3543 1563 3544
rect 1557 3539 1559 3543
rect 1579 3540 1580 3544
rect 1575 3539 1580 3540
rect 1582 3543 1589 3544
rect 1582 3539 1585 3543
rect 1604 3541 1606 3544
rect 1600 3539 1606 3541
rect 1608 3543 1613 3544
rect 1608 3539 1609 3543
rect 1968 3573 1973 3574
rect 1972 3569 1973 3573
rect 1975 3573 1981 3574
rect 1975 3569 1977 3573
rect 1994 3573 1999 3574
rect 1998 3569 1999 3573
rect 2001 3573 2007 3574
rect 2001 3569 2003 3573
rect 2023 3570 2024 3574
rect 2019 3569 2024 3570
rect 2026 3573 2033 3574
rect 2026 3569 2029 3573
rect 2048 3571 2050 3574
rect 2044 3569 2050 3571
rect 2052 3573 2057 3574
rect 2052 3569 2053 3573
rect 2145 3574 2150 3575
rect 2149 3570 2150 3574
rect 2152 3574 2158 3575
rect 2152 3570 2154 3574
rect 2171 3574 2176 3575
rect 2175 3570 2176 3574
rect 2178 3574 2184 3575
rect 2178 3570 2180 3574
rect 2200 3571 2201 3575
rect 2196 3570 2201 3571
rect 2203 3574 2210 3575
rect 2203 3570 2206 3574
rect 2225 3572 2227 3575
rect 2221 3570 2227 3572
rect 2229 3574 2234 3575
rect 2229 3570 2230 3574
rect 1377 3449 1378 3452
rect 1373 3447 1378 3449
rect 1380 3450 1387 3452
rect 1380 3447 1382 3450
rect 1386 3447 1387 3450
rect 1389 3449 1391 3452
rect 1389 3447 1395 3449
rect 1419 3449 1420 3452
rect 1415 3447 1420 3449
rect 1422 3448 1425 3452
rect 1422 3447 1429 3448
rect 1693 3462 1694 3465
rect 1563 3455 1564 3458
rect 1559 3453 1564 3455
rect 1566 3456 1573 3458
rect 1566 3453 1568 3456
rect 1572 3453 1573 3456
rect 1575 3455 1577 3458
rect 1575 3453 1581 3455
rect 1689 3460 1694 3462
rect 1696 3460 1704 3465
rect 1706 3463 1724 3465
rect 1706 3460 1712 3463
rect 1605 3455 1606 3458
rect 1601 3453 1606 3455
rect 1608 3454 1611 3458
rect 1608 3453 1615 3454
rect 1716 3460 1724 3463
rect 1998 3480 1999 3483
rect 1994 3478 1999 3480
rect 2001 3481 2008 3483
rect 2001 3478 2003 3481
rect 2007 3478 2008 3481
rect 2010 3480 2012 3483
rect 2010 3478 2016 3480
rect 2040 3480 2041 3483
rect 2036 3478 2041 3480
rect 2043 3479 2046 3483
rect 2043 3478 2050 3479
rect 1749 3462 1750 3465
rect 1745 3460 1750 3462
rect 1752 3461 1755 3465
rect 1752 3460 1759 3461
rect 2314 3493 2315 3496
rect 2184 3486 2185 3489
rect 2180 3484 2185 3486
rect 2187 3487 2194 3489
rect 2187 3484 2189 3487
rect 2193 3484 2194 3487
rect 2196 3486 2198 3489
rect 2196 3484 2202 3486
rect 2310 3491 2315 3493
rect 2317 3491 2325 3496
rect 2327 3494 2345 3496
rect 2327 3491 2333 3494
rect 2226 3486 2227 3489
rect 2222 3484 2227 3486
rect 2229 3485 2232 3489
rect 2229 3484 2236 3485
rect 2337 3491 2345 3494
rect 2370 3493 2371 3496
rect 2366 3491 2371 3493
rect 2373 3492 2376 3496
rect 2373 3491 2380 3492
rect 399 3056 400 3059
rect 395 3054 400 3056
rect 402 3057 409 3059
rect 402 3054 404 3057
rect 408 3054 409 3057
rect 411 3056 413 3059
rect 411 3054 417 3056
rect 441 3056 442 3059
rect 437 3054 442 3056
rect 444 3055 447 3059
rect 444 3054 451 3055
rect 542 3056 543 3059
rect 538 3054 543 3056
rect 545 3057 552 3059
rect 545 3054 547 3057
rect 551 3054 552 3057
rect 554 3056 556 3059
rect 554 3054 560 3056
rect 584 3056 585 3059
rect 580 3054 585 3056
rect 587 3055 590 3059
rect 587 3054 594 3055
rect 705 3056 706 3059
rect 701 3054 706 3056
rect 708 3057 715 3059
rect 708 3054 710 3057
rect 714 3054 715 3057
rect 717 3056 719 3059
rect 717 3054 723 3056
rect 747 3056 748 3059
rect 743 3054 748 3056
rect 750 3055 753 3059
rect 750 3054 757 3055
rect 861 3056 862 3059
rect 857 3054 862 3056
rect 864 3057 871 3059
rect 864 3054 866 3057
rect 870 3054 871 3057
rect 873 3056 875 3059
rect 873 3054 879 3056
rect 903 3056 904 3059
rect 899 3054 904 3056
rect 906 3055 909 3059
rect 906 3054 913 3055
rect 999 3056 1000 3059
rect 995 3054 1000 3056
rect 1002 3057 1009 3059
rect 1002 3054 1004 3057
rect 1008 3054 1009 3057
rect 1011 3056 1013 3059
rect 1011 3054 1017 3056
rect 1041 3056 1042 3059
rect 1037 3054 1042 3056
rect 1044 3055 1047 3059
rect 1044 3054 1051 3055
rect 1142 3056 1143 3059
rect 1138 3054 1143 3056
rect 1145 3057 1152 3059
rect 1145 3054 1147 3057
rect 1151 3054 1152 3057
rect 1154 3056 1156 3059
rect 1154 3054 1160 3056
rect 1184 3056 1185 3059
rect 1180 3054 1185 3056
rect 1187 3055 1190 3059
rect 1187 3054 1194 3055
rect 1305 3056 1306 3059
rect 1301 3054 1306 3056
rect 1308 3057 1315 3059
rect 1308 3054 1310 3057
rect 1314 3054 1315 3057
rect 1317 3056 1319 3059
rect 1317 3054 1323 3056
rect 1347 3056 1348 3059
rect 1343 3054 1348 3056
rect 1350 3055 1353 3059
rect 1350 3054 1357 3055
rect 1461 3056 1462 3059
rect 1457 3054 1462 3056
rect 1464 3057 1471 3059
rect 1464 3054 1466 3057
rect 1470 3054 1471 3057
rect 1473 3056 1475 3059
rect 1473 3054 1479 3056
rect 1503 3056 1504 3059
rect 1499 3054 1504 3056
rect 1506 3055 1509 3059
rect 1506 3054 1513 3055
rect 2965 3249 2970 3250
rect 2969 3245 2970 3249
rect 2972 3249 2978 3250
rect 2972 3245 2974 3249
rect 2991 3249 2996 3250
rect 2995 3245 2996 3249
rect 2998 3249 3004 3250
rect 2998 3245 3000 3249
rect 3020 3246 3021 3250
rect 3016 3245 3021 3246
rect 3023 3249 3030 3250
rect 3023 3245 3026 3249
rect 3045 3247 3047 3250
rect 3041 3245 3047 3247
rect 3049 3249 3054 3250
rect 3049 3245 3050 3249
rect 3142 3250 3147 3251
rect 3146 3246 3147 3250
rect 3149 3250 3155 3251
rect 3149 3246 3151 3250
rect 3168 3250 3173 3251
rect 3172 3246 3173 3250
rect 3175 3250 3181 3251
rect 3175 3246 3177 3250
rect 3197 3247 3198 3251
rect 3193 3246 3198 3247
rect 3200 3250 3207 3251
rect 3200 3246 3203 3250
rect 3222 3248 3224 3251
rect 3218 3246 3224 3248
rect 3226 3250 3231 3251
rect 3226 3246 3227 3250
rect 3528 3256 3533 3257
rect 3532 3252 3533 3256
rect 3535 3256 3541 3257
rect 3535 3252 3537 3256
rect 3554 3256 3559 3257
rect 3558 3252 3559 3256
rect 3561 3256 3567 3257
rect 3561 3252 3563 3256
rect 3583 3253 3584 3257
rect 3579 3252 3584 3253
rect 3586 3256 3593 3257
rect 3586 3252 3589 3256
rect 3608 3254 3610 3257
rect 3604 3252 3610 3254
rect 3612 3256 3617 3257
rect 3612 3252 3613 3256
rect 2995 3156 2996 3159
rect 2991 3154 2996 3156
rect 2998 3157 3005 3159
rect 2998 3154 3000 3157
rect 3004 3154 3005 3157
rect 3007 3156 3009 3159
rect 3007 3154 3013 3156
rect 3037 3156 3038 3159
rect 3033 3154 3038 3156
rect 3040 3155 3043 3159
rect 3040 3154 3047 3155
rect 3705 3257 3710 3258
rect 3709 3253 3710 3257
rect 3712 3257 3718 3258
rect 3712 3253 3714 3257
rect 3731 3257 3736 3258
rect 3735 3253 3736 3257
rect 3738 3257 3744 3258
rect 3738 3253 3740 3257
rect 3760 3254 3761 3258
rect 3756 3253 3761 3254
rect 3763 3257 3770 3258
rect 3763 3253 3766 3257
rect 3785 3255 3787 3258
rect 3781 3253 3787 3255
rect 3789 3257 3794 3258
rect 3789 3253 3790 3257
rect 4104 3242 4109 3243
rect 4108 3238 4109 3242
rect 4111 3242 4117 3243
rect 4111 3238 4113 3242
rect 4130 3242 4135 3243
rect 4134 3238 4135 3242
rect 4137 3242 4143 3243
rect 4137 3238 4139 3242
rect 4159 3239 4160 3243
rect 4155 3238 4160 3239
rect 4162 3242 4169 3243
rect 4162 3238 4165 3242
rect 4184 3240 4186 3243
rect 4180 3238 4186 3240
rect 4188 3242 4193 3243
rect 4188 3238 4189 3242
rect 3311 3169 3312 3172
rect 3181 3162 3182 3165
rect 3177 3160 3182 3162
rect 3184 3163 3191 3165
rect 3184 3160 3186 3163
rect 3190 3160 3191 3163
rect 3193 3162 3195 3165
rect 3193 3160 3199 3162
rect 3307 3167 3312 3169
rect 3314 3167 3322 3172
rect 3324 3170 3342 3172
rect 3324 3167 3330 3170
rect 3223 3162 3224 3165
rect 3219 3160 3224 3162
rect 3226 3161 3229 3165
rect 3226 3160 3233 3161
rect 3334 3167 3342 3170
rect 3367 3169 3368 3172
rect 3363 3167 3368 3169
rect 3370 3168 3373 3172
rect 3370 3167 3377 3168
rect 3558 3163 3559 3166
rect 3554 3161 3559 3163
rect 3561 3164 3568 3166
rect 3561 3161 3563 3164
rect 3567 3161 3568 3164
rect 3570 3163 3572 3166
rect 3570 3161 3576 3163
rect 3600 3163 3601 3166
rect 3596 3161 3601 3163
rect 3603 3162 3606 3166
rect 3603 3161 3610 3162
rect 3874 3176 3875 3179
rect 3744 3169 3745 3172
rect 3740 3167 3745 3169
rect 3747 3170 3754 3172
rect 3747 3167 3749 3170
rect 3753 3167 3754 3170
rect 3756 3169 3758 3172
rect 3756 3167 3762 3169
rect 3870 3174 3875 3176
rect 3877 3174 3885 3179
rect 3887 3177 3905 3179
rect 3887 3174 3893 3177
rect 3786 3169 3787 3172
rect 3782 3167 3787 3169
rect 3789 3168 3792 3172
rect 3789 3167 3796 3168
rect 3897 3174 3905 3177
rect 3930 3176 3931 3179
rect 3926 3174 3931 3176
rect 3933 3175 3936 3179
rect 3933 3174 3940 3175
rect 4281 3243 4286 3244
rect 4285 3239 4286 3243
rect 4288 3243 4294 3244
rect 4288 3239 4290 3243
rect 4307 3243 4312 3244
rect 4311 3239 4312 3243
rect 4314 3243 4320 3244
rect 4314 3239 4316 3243
rect 4336 3240 4337 3244
rect 4332 3239 4337 3240
rect 4339 3243 4346 3244
rect 4339 3239 4342 3243
rect 4361 3241 4363 3244
rect 4357 3239 4363 3241
rect 4365 3243 4370 3244
rect 4365 3239 4366 3243
rect 4725 3273 4730 3274
rect 4729 3269 4730 3273
rect 4732 3273 4738 3274
rect 4732 3269 4734 3273
rect 4751 3273 4756 3274
rect 4755 3269 4756 3273
rect 4758 3273 4764 3274
rect 4758 3269 4760 3273
rect 4780 3270 4781 3274
rect 4776 3269 4781 3270
rect 4783 3273 4790 3274
rect 4783 3269 4786 3273
rect 4805 3271 4807 3274
rect 4801 3269 4807 3271
rect 4809 3273 4814 3274
rect 4809 3269 4810 3273
rect 4902 3274 4907 3275
rect 4906 3270 4907 3274
rect 4909 3274 4915 3275
rect 4909 3270 4911 3274
rect 4928 3274 4933 3275
rect 4932 3270 4933 3274
rect 4935 3274 4941 3275
rect 4935 3270 4937 3274
rect 4957 3271 4958 3275
rect 4953 3270 4958 3271
rect 4960 3274 4967 3275
rect 4960 3270 4963 3274
rect 4982 3272 4984 3275
rect 4978 3270 4984 3272
rect 4986 3274 4991 3275
rect 4986 3270 4987 3274
rect 4134 3149 4135 3152
rect 4130 3147 4135 3149
rect 4137 3150 4144 3152
rect 4137 3147 4139 3150
rect 4143 3147 4144 3150
rect 4146 3149 4148 3152
rect 4146 3147 4152 3149
rect 4176 3149 4177 3152
rect 4172 3147 4177 3149
rect 4179 3148 4182 3152
rect 4179 3147 4186 3148
rect 4450 3162 4451 3165
rect 4320 3155 4321 3158
rect 4316 3153 4321 3155
rect 4323 3156 4330 3158
rect 4323 3153 4325 3156
rect 4329 3153 4330 3156
rect 4332 3155 4334 3158
rect 4332 3153 4338 3155
rect 4446 3160 4451 3162
rect 4453 3160 4461 3165
rect 4463 3163 4481 3165
rect 4463 3160 4469 3163
rect 4362 3155 4363 3158
rect 4358 3153 4363 3155
rect 4365 3154 4368 3158
rect 4365 3153 4372 3154
rect 4473 3160 4481 3163
rect 4755 3180 4756 3183
rect 4751 3178 4756 3180
rect 4758 3181 4765 3183
rect 4758 3178 4760 3181
rect 4764 3178 4765 3181
rect 4767 3180 4769 3183
rect 4767 3178 4773 3180
rect 4797 3180 4798 3183
rect 4793 3178 4798 3180
rect 4800 3179 4803 3183
rect 4800 3178 4807 3179
rect 4506 3162 4507 3165
rect 4502 3160 4507 3162
rect 4509 3161 4512 3165
rect 4509 3160 4516 3161
rect 5071 3193 5072 3196
rect 4941 3186 4942 3189
rect 4937 3184 4942 3186
rect 4944 3187 4951 3189
rect 4944 3184 4946 3187
rect 4950 3184 4951 3187
rect 4953 3186 4955 3189
rect 4953 3184 4959 3186
rect 5067 3191 5072 3193
rect 5074 3191 5082 3196
rect 5084 3194 5102 3196
rect 5084 3191 5090 3194
rect 4983 3186 4984 3189
rect 4979 3184 4984 3186
rect 4986 3185 4989 3189
rect 4986 3184 4993 3185
rect 5094 3191 5102 3194
rect 5127 3193 5128 3196
rect 5123 3191 5128 3193
rect 5130 3192 5133 3196
rect 5130 3191 5137 3192
rect 241 2988 242 2991
rect 237 2986 242 2988
rect 244 2989 251 2991
rect 244 2986 246 2989
rect 250 2986 251 2989
rect 253 2988 255 2991
rect 253 2986 259 2988
rect 283 2988 284 2991
rect 279 2986 284 2988
rect 286 2987 289 2991
rect 286 2986 293 2987
rect 193 2934 194 2938
rect 196 2934 197 2938
rect 104 2904 105 2907
rect 100 2902 105 2904
rect 107 2905 114 2907
rect 107 2902 109 2905
rect 113 2902 114 2905
rect 116 2904 118 2907
rect 116 2902 122 2904
rect 146 2904 147 2907
rect 142 2902 147 2904
rect 149 2903 152 2907
rect 149 2902 156 2903
rect 240 2907 241 2910
rect 236 2905 241 2907
rect 243 2908 250 2910
rect 243 2905 245 2908
rect 249 2905 250 2908
rect 252 2907 254 2910
rect 252 2905 258 2907
rect 282 2907 283 2910
rect 278 2905 283 2907
rect 285 2906 288 2910
rect 285 2905 292 2906
rect 193 2851 194 2855
rect 196 2851 197 2855
rect 399 2914 400 2917
rect 395 2912 400 2914
rect 402 2915 409 2917
rect 402 2912 404 2915
rect 408 2912 409 2915
rect 411 2914 413 2917
rect 411 2912 417 2914
rect 441 2914 442 2917
rect 437 2912 442 2914
rect 444 2913 447 2917
rect 444 2912 451 2913
rect 542 2914 543 2917
rect 538 2912 543 2914
rect 545 2915 552 2917
rect 545 2912 547 2915
rect 551 2912 552 2915
rect 554 2914 556 2917
rect 554 2912 560 2914
rect 584 2914 585 2917
rect 580 2912 585 2914
rect 587 2913 590 2917
rect 587 2912 594 2913
rect 705 2914 706 2917
rect 701 2912 706 2914
rect 708 2915 715 2917
rect 708 2912 710 2915
rect 714 2912 715 2915
rect 717 2914 719 2917
rect 717 2912 723 2914
rect 747 2914 748 2917
rect 743 2912 748 2914
rect 750 2913 753 2917
rect 750 2912 757 2913
rect 861 2914 862 2917
rect 857 2912 862 2914
rect 864 2915 871 2917
rect 864 2912 866 2915
rect 870 2912 871 2915
rect 873 2914 875 2917
rect 873 2912 879 2914
rect 903 2914 904 2917
rect 899 2912 904 2914
rect 906 2913 909 2917
rect 906 2912 913 2913
rect 999 2914 1000 2917
rect 995 2912 1000 2914
rect 1002 2915 1009 2917
rect 1002 2912 1004 2915
rect 1008 2912 1009 2915
rect 1011 2914 1013 2917
rect 1011 2912 1017 2914
rect 1041 2914 1042 2917
rect 1037 2912 1042 2914
rect 1044 2913 1047 2917
rect 1044 2912 1051 2913
rect 1142 2914 1143 2917
rect 1138 2912 1143 2914
rect 1145 2915 1152 2917
rect 1145 2912 1147 2915
rect 1151 2912 1152 2915
rect 1154 2914 1156 2917
rect 1154 2912 1160 2914
rect 1184 2914 1185 2917
rect 1180 2912 1185 2914
rect 1187 2913 1190 2917
rect 1187 2912 1194 2913
rect 1305 2914 1306 2917
rect 1301 2912 1306 2914
rect 1308 2915 1315 2917
rect 1308 2912 1310 2915
rect 1314 2912 1315 2915
rect 1317 2914 1319 2917
rect 1317 2912 1323 2914
rect 1347 2914 1348 2917
rect 1343 2912 1348 2914
rect 1350 2913 1353 2917
rect 1350 2912 1357 2913
rect 1461 2914 1462 2917
rect 1457 2912 1462 2914
rect 1464 2915 1471 2917
rect 1464 2912 1466 2915
rect 1470 2912 1471 2915
rect 1473 2914 1475 2917
rect 1473 2912 1479 2914
rect 1503 2914 1504 2917
rect 1499 2912 1504 2914
rect 1506 2913 1509 2917
rect 1506 2912 1513 2913
rect 1692 2939 1697 2940
rect 1696 2935 1697 2939
rect 1699 2939 1705 2940
rect 1699 2935 1701 2939
rect 1718 2939 1723 2940
rect 1722 2935 1723 2939
rect 1725 2939 1731 2940
rect 1725 2935 1727 2939
rect 1747 2936 1748 2940
rect 1743 2935 1748 2936
rect 1750 2939 1757 2940
rect 1750 2935 1753 2939
rect 1772 2937 1774 2940
rect 1768 2935 1774 2937
rect 1776 2939 1781 2940
rect 1776 2935 1777 2939
rect 1887 2940 1892 2941
rect 1891 2936 1892 2940
rect 1894 2940 1900 2941
rect 1894 2936 1896 2940
rect 1913 2940 1918 2941
rect 1917 2936 1918 2940
rect 1920 2940 1926 2941
rect 1920 2936 1922 2940
rect 1942 2937 1943 2941
rect 1938 2936 1943 2937
rect 1945 2940 1952 2941
rect 1945 2936 1948 2940
rect 1967 2938 1969 2941
rect 1963 2936 1969 2938
rect 1971 2940 1976 2941
rect 1971 2936 1972 2940
rect 2100 2939 2105 2940
rect 2104 2935 2105 2939
rect 2107 2939 2113 2940
rect 2107 2935 2109 2939
rect 2126 2939 2131 2940
rect 2130 2935 2131 2939
rect 2133 2939 2139 2940
rect 2133 2935 2135 2939
rect 2155 2936 2156 2940
rect 2151 2935 2156 2936
rect 2158 2939 2165 2940
rect 2158 2935 2161 2939
rect 2180 2937 2182 2940
rect 2176 2935 2182 2937
rect 2184 2939 2189 2940
rect 2184 2935 2185 2939
rect 2301 2940 2306 2941
rect 2305 2936 2306 2940
rect 2308 2940 2314 2941
rect 2308 2936 2310 2940
rect 2327 2940 2332 2941
rect 2331 2936 2332 2940
rect 2334 2940 2340 2941
rect 2334 2936 2336 2940
rect 2356 2937 2357 2941
rect 2352 2936 2357 2937
rect 2359 2940 2366 2941
rect 2359 2936 2362 2940
rect 2381 2938 2383 2941
rect 2377 2936 2383 2938
rect 2385 2940 2390 2941
rect 2385 2936 2386 2940
rect 244 2816 245 2819
rect 240 2814 245 2816
rect 247 2817 254 2819
rect 247 2814 249 2817
rect 253 2814 254 2817
rect 256 2816 258 2819
rect 256 2814 262 2816
rect 286 2816 287 2819
rect 282 2814 287 2816
rect 289 2815 292 2819
rect 289 2814 296 2815
rect 399 2765 400 2768
rect 395 2763 400 2765
rect 402 2766 409 2768
rect 402 2763 404 2766
rect 408 2763 409 2766
rect 411 2765 413 2768
rect 411 2763 417 2765
rect 441 2765 442 2768
rect 437 2763 442 2765
rect 444 2764 447 2768
rect 444 2763 451 2764
rect 542 2765 543 2768
rect 538 2763 543 2765
rect 545 2766 552 2768
rect 545 2763 547 2766
rect 551 2763 552 2766
rect 554 2765 556 2768
rect 554 2763 560 2765
rect 584 2765 585 2768
rect 580 2763 585 2765
rect 587 2764 590 2768
rect 587 2763 594 2764
rect 705 2765 706 2768
rect 701 2763 706 2765
rect 708 2766 715 2768
rect 708 2763 710 2766
rect 714 2763 715 2766
rect 717 2765 719 2768
rect 717 2763 723 2765
rect 747 2765 748 2768
rect 743 2763 748 2765
rect 750 2764 753 2768
rect 750 2763 757 2764
rect 861 2765 862 2768
rect 857 2763 862 2765
rect 864 2766 871 2768
rect 864 2763 866 2766
rect 870 2763 871 2766
rect 873 2765 875 2768
rect 873 2763 879 2765
rect 903 2765 904 2768
rect 899 2763 904 2765
rect 906 2764 909 2768
rect 906 2763 913 2764
rect 999 2765 1000 2768
rect 995 2763 1000 2765
rect 1002 2766 1009 2768
rect 1002 2763 1004 2766
rect 1008 2763 1009 2766
rect 1011 2765 1013 2768
rect 1011 2763 1017 2765
rect 1041 2765 1042 2768
rect 1037 2763 1042 2765
rect 1044 2764 1047 2768
rect 1044 2763 1051 2764
rect 1142 2765 1143 2768
rect 1138 2763 1143 2765
rect 1145 2766 1152 2768
rect 1145 2763 1147 2766
rect 1151 2763 1152 2766
rect 1154 2765 1156 2768
rect 1154 2763 1160 2765
rect 1184 2765 1185 2768
rect 1180 2763 1185 2765
rect 1187 2764 1190 2768
rect 1187 2763 1194 2764
rect 1305 2765 1306 2768
rect 1301 2763 1306 2765
rect 1308 2766 1315 2768
rect 1308 2763 1310 2766
rect 1314 2763 1315 2766
rect 1317 2765 1319 2768
rect 1317 2763 1323 2765
rect 1347 2765 1348 2768
rect 1343 2763 1348 2765
rect 1350 2764 1353 2768
rect 1350 2763 1357 2764
rect 1461 2765 1462 2768
rect 1457 2763 1462 2765
rect 1464 2766 1471 2768
rect 1464 2763 1466 2766
rect 1470 2763 1471 2766
rect 1473 2765 1475 2768
rect 1473 2763 1479 2765
rect 1503 2765 1504 2768
rect 1499 2763 1504 2765
rect 1506 2764 1509 2768
rect 1506 2763 1513 2764
rect 2360 2746 2369 2752
rect 2364 2742 2369 2746
rect 2371 2746 2384 2752
rect 2371 2742 2373 2746
rect 2377 2742 2384 2746
rect 2386 2746 2399 2752
rect 2386 2742 2390 2746
rect 2394 2742 2399 2746
rect 2401 2746 2414 2752
rect 2401 2742 2405 2746
rect 2409 2742 2414 2746
rect 2416 2746 2428 2752
rect 2416 2742 2420 2746
rect 2424 2742 2428 2746
rect 2430 2746 2439 2752
rect 2430 2742 2435 2746
rect 2445 2746 2454 2752
rect 2449 2742 2454 2746
rect 2456 2746 2465 2752
rect 2456 2742 2461 2746
rect 2122 2688 2123 2692
rect 2125 2688 2126 2692
rect 399 2640 400 2643
rect 395 2638 400 2640
rect 402 2641 409 2643
rect 402 2638 404 2641
rect 408 2638 409 2641
rect 411 2640 413 2643
rect 411 2638 417 2640
rect 441 2640 442 2643
rect 437 2638 442 2640
rect 444 2639 447 2643
rect 444 2638 451 2639
rect 542 2640 543 2643
rect 538 2638 543 2640
rect 545 2641 552 2643
rect 545 2638 547 2641
rect 551 2638 552 2641
rect 554 2640 556 2643
rect 554 2638 560 2640
rect 584 2640 585 2643
rect 580 2638 585 2640
rect 587 2639 590 2643
rect 587 2638 594 2639
rect 705 2640 706 2643
rect 701 2638 706 2640
rect 708 2641 715 2643
rect 708 2638 710 2641
rect 714 2638 715 2641
rect 717 2640 719 2643
rect 717 2638 723 2640
rect 747 2640 748 2643
rect 743 2638 748 2640
rect 750 2639 753 2643
rect 750 2638 757 2639
rect 861 2640 862 2643
rect 857 2638 862 2640
rect 864 2641 871 2643
rect 864 2638 866 2641
rect 870 2638 871 2641
rect 873 2640 875 2643
rect 873 2638 879 2640
rect 903 2640 904 2643
rect 899 2638 904 2640
rect 906 2639 909 2643
rect 906 2638 913 2639
rect 999 2640 1000 2643
rect 995 2638 1000 2640
rect 1002 2641 1009 2643
rect 1002 2638 1004 2641
rect 1008 2638 1009 2641
rect 1011 2640 1013 2643
rect 1011 2638 1017 2640
rect 1041 2640 1042 2643
rect 1037 2638 1042 2640
rect 1044 2639 1047 2643
rect 1044 2638 1051 2639
rect 1142 2640 1143 2643
rect 1138 2638 1143 2640
rect 1145 2641 1152 2643
rect 1145 2638 1147 2641
rect 1151 2638 1152 2641
rect 1154 2640 1156 2643
rect 1154 2638 1160 2640
rect 1184 2640 1185 2643
rect 1180 2638 1185 2640
rect 1187 2639 1190 2643
rect 1187 2638 1194 2639
rect 1305 2640 1306 2643
rect 1301 2638 1306 2640
rect 1308 2641 1315 2643
rect 1308 2638 1310 2641
rect 1314 2638 1315 2641
rect 1317 2640 1319 2643
rect 1317 2638 1323 2640
rect 1347 2640 1348 2643
rect 1343 2638 1348 2640
rect 1350 2639 1353 2643
rect 1350 2638 1357 2639
rect 1461 2640 1462 2643
rect 1457 2638 1462 2640
rect 1464 2641 1471 2643
rect 1464 2638 1466 2641
rect 1470 2638 1471 2641
rect 1473 2640 1475 2643
rect 1473 2638 1479 2640
rect 1503 2640 1504 2643
rect 1499 2638 1504 2640
rect 1506 2639 1509 2643
rect 1506 2638 1513 2639
rect 781 2281 782 2284
rect 777 2279 782 2281
rect 784 2282 791 2284
rect 784 2279 786 2282
rect 790 2279 791 2282
rect 793 2281 795 2284
rect 793 2279 799 2281
rect 823 2281 824 2284
rect 819 2279 824 2281
rect 826 2280 829 2284
rect 826 2279 833 2280
rect 924 2281 925 2284
rect 920 2279 925 2281
rect 927 2282 934 2284
rect 927 2279 929 2282
rect 933 2279 934 2282
rect 936 2281 938 2284
rect 936 2279 942 2281
rect 966 2281 967 2284
rect 962 2279 967 2281
rect 969 2280 972 2284
rect 969 2279 976 2280
rect 1087 2281 1088 2284
rect 1083 2279 1088 2281
rect 1090 2282 1097 2284
rect 1090 2279 1092 2282
rect 1096 2279 1097 2282
rect 1099 2281 1101 2284
rect 1099 2279 1105 2281
rect 1129 2281 1130 2284
rect 1125 2279 1130 2281
rect 1132 2280 1135 2284
rect 1132 2279 1139 2280
rect 1243 2281 1244 2284
rect 1239 2279 1244 2281
rect 1246 2282 1253 2284
rect 1246 2279 1248 2282
rect 1252 2279 1253 2282
rect 1255 2281 1257 2284
rect 1255 2279 1261 2281
rect 1285 2281 1286 2284
rect 1281 2279 1286 2281
rect 1288 2280 1291 2284
rect 1288 2279 1295 2280
rect 2491 2646 2500 2652
rect 2495 2642 2500 2646
rect 2502 2646 2515 2652
rect 2502 2642 2506 2646
rect 2511 2642 2515 2646
rect 2517 2646 2535 2652
rect 2517 2642 2524 2646
rect 2528 2642 2535 2646
rect 2537 2646 2545 2652
rect 2537 2642 2539 2646
rect 2543 2642 2545 2646
rect 2547 2646 2557 2652
rect 2547 2642 2553 2646
rect 2562 2646 2571 2652
rect 2566 2642 2571 2646
rect 2573 2646 2582 2652
rect 2573 2642 2578 2646
rect 2810 2696 2818 2699
rect 2814 2692 2818 2696
rect 2820 2692 2830 2699
rect 2832 2692 2845 2699
rect 2847 2692 2855 2699
rect 2857 2696 2866 2699
rect 2857 2692 2862 2696
rect 2870 2696 2878 2699
rect 2874 2692 2878 2696
rect 2880 2696 2887 2699
rect 2880 2692 2883 2696
rect 2124 2622 2125 2626
rect 2127 2622 2128 2626
rect 2629 2608 2638 2614
rect 2127 2555 2128 2559
rect 2130 2555 2131 2559
rect 2127 2488 2128 2492
rect 2130 2488 2131 2492
rect 2145 2383 2146 2387
rect 2148 2383 2149 2387
rect 2041 2350 2046 2351
rect 2045 2346 2046 2350
rect 2048 2350 2054 2351
rect 2048 2346 2050 2350
rect 2060 2350 2065 2351
rect 2064 2346 2065 2350
rect 2067 2350 2073 2351
rect 2067 2346 2069 2350
rect 2085 2350 2090 2351
rect 2089 2346 2090 2350
rect 2092 2350 2098 2351
rect 2092 2346 2094 2350
rect 2104 2350 2109 2351
rect 2108 2346 2109 2350
rect 2111 2350 2117 2351
rect 2111 2346 2113 2350
rect 2147 2222 2148 2226
rect 2150 2222 2151 2226
rect 2043 2189 2048 2190
rect 2047 2185 2048 2189
rect 2050 2189 2056 2190
rect 2050 2185 2052 2189
rect 2062 2189 2067 2190
rect 2066 2185 2067 2189
rect 2069 2189 2075 2190
rect 2069 2185 2071 2189
rect 2087 2189 2092 2190
rect 2091 2185 2092 2189
rect 2094 2189 2100 2190
rect 2094 2185 2096 2189
rect 2106 2189 2111 2190
rect 2110 2185 2111 2189
rect 2113 2189 2119 2190
rect 2113 2185 2115 2189
rect 2633 2604 2638 2608
rect 2640 2608 2653 2614
rect 2640 2604 2644 2608
rect 2649 2604 2653 2608
rect 2655 2608 2673 2614
rect 2655 2604 2662 2608
rect 2666 2604 2673 2608
rect 2675 2608 2683 2614
rect 2675 2604 2679 2608
rect 2688 2608 2697 2614
rect 2692 2604 2697 2608
rect 2699 2608 2708 2614
rect 2699 2604 2704 2608
rect 2758 2568 2764 2569
rect 2762 2564 2764 2568
rect 2766 2565 2769 2569
rect 2766 2564 2773 2565
rect 2779 2568 2785 2569
rect 2783 2564 2785 2568
rect 2787 2565 2790 2569
rect 2810 2565 2811 2569
rect 2813 2565 2814 2569
rect 2787 2564 2794 2565
rect 2738 2172 2747 2178
rect 2742 2168 2747 2172
rect 2749 2172 2762 2178
rect 2749 2168 2753 2172
rect 2758 2168 2762 2172
rect 2764 2172 2782 2178
rect 2764 2168 2771 2172
rect 2775 2168 2782 2172
rect 2784 2172 2792 2178
rect 2784 2168 2786 2172
rect 2790 2168 2792 2172
rect 2794 2172 2804 2178
rect 2794 2168 2800 2172
rect 2809 2172 2818 2178
rect 2813 2168 2818 2172
rect 2820 2172 2829 2178
rect 2820 2168 2825 2172
rect 2905 2166 2906 2169
rect 2901 2164 2906 2166
rect 2908 2167 2917 2169
rect 2908 2164 2912 2167
rect 2916 2164 2917 2167
rect 2919 2166 2921 2169
rect 2919 2164 2925 2166
rect 2947 2166 2948 2169
rect 2943 2164 2948 2166
rect 2950 2165 2953 2169
rect 2950 2164 2957 2165
rect 2146 2068 2147 2072
rect 2149 2068 2150 2072
rect 2042 2035 2047 2036
rect 2046 2031 2047 2035
rect 2049 2035 2055 2036
rect 2049 2031 2051 2035
rect 2061 2035 2066 2036
rect 2065 2031 2066 2035
rect 2068 2035 2074 2036
rect 2068 2031 2070 2035
rect 2086 2035 2091 2036
rect 2090 2031 2091 2035
rect 2093 2035 2099 2036
rect 2093 2031 2095 2035
rect 2105 2035 2110 2036
rect 2109 2031 2110 2035
rect 2112 2035 2118 2036
rect 2112 2031 2114 2035
rect 2146 1920 2147 1924
rect 2149 1920 2150 1924
rect 2801 1916 2809 1919
rect 2805 1912 2809 1916
rect 2811 1912 2821 1919
rect 2823 1912 2836 1919
rect 2838 1912 2846 1919
rect 2848 1916 2857 1919
rect 2848 1912 2853 1916
rect 2861 1916 2869 1919
rect 2865 1912 2869 1916
rect 2871 1916 2878 1919
rect 2871 1912 2874 1916
rect 2042 1887 2047 1888
rect 2046 1883 2047 1887
rect 2049 1887 2055 1888
rect 2049 1883 2051 1887
rect 2061 1887 2066 1888
rect 2065 1883 2066 1887
rect 2068 1887 2074 1888
rect 2068 1883 2070 1887
rect 2086 1887 2091 1888
rect 2090 1883 2091 1887
rect 2093 1887 2099 1888
rect 2093 1883 2095 1887
rect 2105 1887 2110 1888
rect 2109 1883 2110 1887
rect 2112 1887 2118 1888
rect 2112 1883 2114 1887
rect 2575 1857 2584 1863
rect 2579 1853 2584 1857
rect 2586 1857 2599 1863
rect 2586 1853 2588 1857
rect 2592 1853 2599 1857
rect 2601 1857 2614 1863
rect 2601 1853 2605 1857
rect 2609 1853 2614 1857
rect 2616 1857 2629 1863
rect 2616 1853 2620 1857
rect 2624 1853 2629 1857
rect 2631 1857 2643 1863
rect 2631 1853 2635 1857
rect 2639 1853 2643 1857
rect 2645 1857 2654 1863
rect 2645 1853 2650 1857
rect 2660 1857 2669 1863
rect 2664 1853 2669 1857
rect 2671 1857 2680 1863
rect 2671 1853 2676 1857
rect 2122 1793 2123 1797
rect 2125 1793 2126 1797
rect 2443 1773 2452 1779
rect 2447 1769 2452 1773
rect 2454 1773 2467 1779
rect 2454 1769 2458 1773
rect 2463 1769 2467 1773
rect 2469 1773 2487 1779
rect 2469 1769 2476 1773
rect 2480 1769 2487 1773
rect 2489 1773 2497 1779
rect 2489 1769 2491 1773
rect 2495 1769 2497 1773
rect 2499 1773 2509 1779
rect 2499 1769 2505 1773
rect 2514 1773 2523 1779
rect 2518 1769 2523 1773
rect 2525 1773 2534 1779
rect 2525 1769 2530 1773
rect 2124 1727 2125 1731
rect 2127 1727 2128 1731
rect 2302 1698 2311 1704
rect 2306 1694 2311 1698
rect 2313 1698 2326 1704
rect 2313 1694 2317 1698
rect 2322 1694 2326 1698
rect 2328 1698 2346 1704
rect 2328 1694 2335 1698
rect 2339 1694 2346 1698
rect 2348 1698 2356 1704
rect 2348 1694 2352 1698
rect 2361 1698 2370 1704
rect 2365 1694 2370 1698
rect 2372 1698 2381 1704
rect 2372 1694 2377 1698
rect 2127 1660 2128 1664
rect 2130 1660 2131 1664
rect 2207 1624 2213 1625
rect 2211 1620 2213 1624
rect 2215 1621 2218 1625
rect 2215 1620 2222 1621
rect 2228 1624 2234 1625
rect 2232 1620 2234 1624
rect 2236 1621 2239 1625
rect 2259 1621 2260 1625
rect 2262 1621 2263 1625
rect 2236 1620 2243 1621
rect 2127 1593 2128 1597
rect 2130 1593 2131 1597
<< ndcontact >>
rect 208 3515 212 3519
rect 217 3515 221 3519
rect 234 3515 238 3519
rect 243 3515 247 3519
rect 259 3514 263 3518
rect 269 3515 273 3519
rect 284 3514 288 3518
rect 293 3515 297 3519
rect 385 3516 389 3520
rect 394 3516 398 3520
rect 411 3516 415 3520
rect 420 3516 424 3520
rect 436 3515 440 3519
rect 446 3516 450 3520
rect 461 3515 465 3519
rect 470 3516 474 3520
rect 771 3522 775 3526
rect 780 3522 784 3526
rect 797 3522 801 3526
rect 806 3522 810 3526
rect 822 3521 826 3525
rect 832 3522 836 3526
rect 847 3521 851 3525
rect 856 3522 860 3526
rect 948 3523 952 3527
rect 957 3523 961 3527
rect 974 3523 978 3527
rect 983 3523 987 3527
rect 999 3522 1003 3526
rect 1009 3523 1013 3527
rect 1024 3522 1028 3526
rect 1033 3523 1037 3527
rect 1347 3508 1351 3512
rect 1356 3508 1360 3512
rect 1373 3508 1377 3512
rect 1382 3508 1386 3512
rect 1398 3507 1402 3511
rect 1408 3508 1412 3512
rect 1423 3507 1427 3511
rect 1432 3508 1436 3512
rect 420 3429 424 3433
rect 438 3430 442 3434
rect 234 3423 238 3427
rect 252 3424 256 3428
rect 276 3422 280 3426
rect 286 3425 290 3429
rect 462 3428 466 3432
rect 472 3431 476 3435
rect 550 3428 554 3432
rect 560 3430 564 3434
rect 983 3436 987 3440
rect 1001 3437 1005 3441
rect 573 3429 577 3433
rect 606 3427 610 3431
rect 616 3430 620 3434
rect 797 3430 801 3434
rect 815 3431 819 3435
rect 839 3429 843 3433
rect 849 3432 853 3436
rect 1025 3435 1029 3439
rect 1035 3438 1039 3442
rect 1113 3435 1117 3439
rect 1123 3437 1127 3441
rect 1524 3509 1528 3513
rect 1533 3509 1537 3513
rect 1550 3509 1554 3513
rect 1559 3509 1563 3513
rect 1575 3508 1579 3512
rect 1585 3509 1589 3513
rect 1600 3508 1604 3512
rect 1609 3509 1613 3513
rect 1968 3539 1972 3543
rect 1977 3539 1981 3543
rect 1994 3539 1998 3543
rect 2003 3539 2007 3543
rect 2019 3538 2023 3542
rect 2029 3539 2033 3543
rect 2044 3538 2048 3542
rect 2053 3539 2057 3543
rect 2145 3540 2149 3544
rect 2154 3540 2158 3544
rect 2171 3540 2175 3544
rect 2180 3540 2184 3544
rect 2196 3539 2200 3543
rect 2206 3540 2210 3544
rect 2221 3539 2225 3543
rect 2230 3540 2234 3544
rect 1136 3436 1140 3440
rect 1169 3434 1173 3438
rect 1179 3437 1183 3441
rect 1559 3422 1563 3426
rect 1577 3423 1581 3427
rect 1373 3416 1377 3420
rect 1391 3417 1395 3421
rect 1415 3415 1419 3419
rect 1425 3418 1429 3422
rect 1601 3421 1605 3425
rect 1611 3424 1615 3428
rect 1689 3421 1693 3425
rect 1699 3423 1703 3427
rect 2180 3453 2184 3457
rect 2198 3454 2202 3458
rect 1994 3447 1998 3451
rect 2012 3448 2016 3452
rect 2036 3446 2040 3450
rect 2046 3449 2050 3453
rect 2222 3452 2226 3456
rect 2232 3455 2236 3459
rect 1712 3422 1716 3426
rect 1745 3420 1749 3424
rect 1755 3423 1759 3427
rect 2310 3452 2314 3456
rect 2320 3454 2324 3458
rect 2333 3453 2337 3457
rect 2366 3451 2370 3455
rect 2376 3454 2380 3458
rect 395 3023 399 3027
rect 413 3024 417 3028
rect 437 3022 441 3026
rect 447 3025 451 3029
rect 538 3023 542 3027
rect 556 3024 560 3028
rect 580 3022 584 3026
rect 590 3025 594 3029
rect 701 3023 705 3027
rect 719 3024 723 3028
rect 743 3022 747 3026
rect 753 3025 757 3029
rect 857 3023 861 3027
rect 875 3024 879 3028
rect 899 3022 903 3026
rect 909 3025 913 3029
rect 995 3023 999 3027
rect 1013 3024 1017 3028
rect 1037 3022 1041 3026
rect 1047 3025 1051 3029
rect 1138 3023 1142 3027
rect 1156 3024 1160 3028
rect 1180 3022 1184 3026
rect 1190 3025 1194 3029
rect 1301 3023 1305 3027
rect 1319 3024 1323 3028
rect 1343 3022 1347 3026
rect 1353 3025 1357 3029
rect 1457 3023 1461 3027
rect 1475 3024 1479 3028
rect 1499 3022 1503 3026
rect 1509 3025 1513 3029
rect 2965 3215 2969 3219
rect 2974 3215 2978 3219
rect 2991 3215 2995 3219
rect 3000 3215 3004 3219
rect 3016 3214 3020 3218
rect 3026 3215 3030 3219
rect 3041 3214 3045 3218
rect 3050 3215 3054 3219
rect 3142 3216 3146 3220
rect 3151 3216 3155 3220
rect 3168 3216 3172 3220
rect 3177 3216 3181 3220
rect 3193 3215 3197 3219
rect 3203 3216 3207 3220
rect 3218 3215 3222 3219
rect 3227 3216 3231 3220
rect 3528 3222 3532 3226
rect 3537 3222 3541 3226
rect 3554 3222 3558 3226
rect 3563 3222 3567 3226
rect 3579 3221 3583 3225
rect 3589 3222 3593 3226
rect 3604 3221 3608 3225
rect 3613 3222 3617 3226
rect 3705 3223 3709 3227
rect 3714 3223 3718 3227
rect 3731 3223 3735 3227
rect 3740 3223 3744 3227
rect 3756 3222 3760 3226
rect 3766 3223 3770 3227
rect 3781 3222 3785 3226
rect 3790 3223 3794 3227
rect 4104 3208 4108 3212
rect 4113 3208 4117 3212
rect 4130 3208 4134 3212
rect 4139 3208 4143 3212
rect 4155 3207 4159 3211
rect 4165 3208 4169 3212
rect 4180 3207 4184 3211
rect 4189 3208 4193 3212
rect 3177 3129 3181 3133
rect 3195 3130 3199 3134
rect 2991 3123 2995 3127
rect 3009 3124 3013 3128
rect 3033 3122 3037 3126
rect 3043 3125 3047 3129
rect 3219 3128 3223 3132
rect 3229 3131 3233 3135
rect 3307 3128 3311 3132
rect 3317 3130 3321 3134
rect 3740 3136 3744 3140
rect 3758 3137 3762 3141
rect 3330 3129 3334 3133
rect 3363 3127 3367 3131
rect 3373 3130 3377 3134
rect 3554 3130 3558 3134
rect 3572 3131 3576 3135
rect 3596 3129 3600 3133
rect 3606 3132 3610 3136
rect 3782 3135 3786 3139
rect 3792 3138 3796 3142
rect 3870 3135 3874 3139
rect 3880 3137 3884 3141
rect 4281 3209 4285 3213
rect 4290 3209 4294 3213
rect 4307 3209 4311 3213
rect 4316 3209 4320 3213
rect 4332 3208 4336 3212
rect 4342 3209 4346 3213
rect 4357 3208 4361 3212
rect 4366 3209 4370 3213
rect 4725 3239 4729 3243
rect 4734 3239 4738 3243
rect 4751 3239 4755 3243
rect 4760 3239 4764 3243
rect 4776 3238 4780 3242
rect 4786 3239 4790 3243
rect 4801 3238 4805 3242
rect 4810 3239 4814 3243
rect 4902 3240 4906 3244
rect 4911 3240 4915 3244
rect 4928 3240 4932 3244
rect 4937 3240 4941 3244
rect 4953 3239 4957 3243
rect 4963 3240 4967 3244
rect 4978 3239 4982 3243
rect 4987 3240 4991 3244
rect 3893 3136 3897 3140
rect 3926 3134 3930 3138
rect 3936 3137 3940 3141
rect 4316 3122 4320 3126
rect 4334 3123 4338 3127
rect 4130 3116 4134 3120
rect 4148 3117 4152 3121
rect 4172 3115 4176 3119
rect 4182 3118 4186 3122
rect 4358 3121 4362 3125
rect 4368 3124 4372 3128
rect 4446 3121 4450 3125
rect 4456 3123 4460 3127
rect 4937 3153 4941 3157
rect 4955 3154 4959 3158
rect 4751 3147 4755 3151
rect 4769 3148 4773 3152
rect 4793 3146 4797 3150
rect 4803 3149 4807 3153
rect 4979 3152 4983 3156
rect 4989 3155 4993 3159
rect 4469 3122 4473 3126
rect 4502 3120 4506 3124
rect 4512 3123 4516 3127
rect 5067 3152 5071 3156
rect 5077 3154 5081 3158
rect 5090 3153 5094 3157
rect 5123 3151 5127 3155
rect 5133 3154 5137 3158
rect 237 2955 241 2959
rect 255 2956 259 2960
rect 279 2954 283 2958
rect 289 2957 293 2961
rect 100 2871 104 2875
rect 118 2872 122 2876
rect 142 2870 146 2874
rect 152 2873 156 2877
rect 189 2911 193 2915
rect 197 2911 201 2915
rect 236 2874 240 2878
rect 254 2875 258 2879
rect 278 2873 282 2877
rect 288 2876 292 2880
rect 395 2881 399 2885
rect 413 2882 417 2886
rect 437 2880 441 2884
rect 447 2883 451 2887
rect 538 2881 542 2885
rect 556 2882 560 2886
rect 580 2880 584 2884
rect 590 2883 594 2887
rect 701 2881 705 2885
rect 719 2882 723 2886
rect 743 2880 747 2884
rect 753 2883 757 2887
rect 857 2881 861 2885
rect 875 2882 879 2886
rect 899 2880 903 2884
rect 909 2883 913 2887
rect 995 2881 999 2885
rect 1013 2882 1017 2886
rect 1037 2880 1041 2884
rect 1047 2883 1051 2887
rect 1138 2881 1142 2885
rect 1156 2882 1160 2886
rect 1180 2880 1184 2884
rect 1190 2883 1194 2887
rect 1301 2881 1305 2885
rect 1319 2882 1323 2886
rect 1343 2880 1347 2884
rect 1353 2883 1357 2887
rect 1457 2881 1461 2885
rect 1475 2882 1479 2886
rect 1499 2880 1503 2884
rect 1509 2883 1513 2887
rect 1692 2905 1696 2909
rect 1701 2905 1705 2909
rect 1718 2905 1722 2909
rect 1727 2905 1731 2909
rect 1743 2904 1747 2908
rect 1753 2905 1757 2909
rect 1768 2904 1772 2908
rect 1777 2905 1781 2909
rect 1887 2906 1891 2910
rect 1896 2906 1900 2910
rect 1913 2906 1917 2910
rect 1922 2906 1926 2910
rect 1938 2905 1942 2909
rect 1948 2906 1952 2910
rect 1963 2905 1967 2909
rect 1972 2906 1976 2910
rect 2100 2905 2104 2909
rect 2109 2905 2113 2909
rect 2126 2905 2130 2909
rect 2135 2905 2139 2909
rect 2151 2904 2155 2908
rect 2161 2905 2165 2909
rect 2176 2904 2180 2908
rect 2185 2905 2189 2909
rect 2301 2906 2305 2910
rect 2310 2906 2314 2910
rect 2327 2906 2331 2910
rect 2336 2906 2340 2910
rect 2352 2905 2356 2909
rect 2362 2906 2366 2910
rect 2377 2905 2381 2909
rect 2386 2906 2390 2910
rect 189 2829 193 2833
rect 197 2829 201 2833
rect 240 2783 244 2787
rect 258 2784 262 2788
rect 282 2782 286 2786
rect 292 2785 296 2789
rect 395 2732 399 2736
rect 413 2733 417 2737
rect 437 2731 441 2735
rect 447 2734 451 2738
rect 538 2732 542 2736
rect 556 2733 560 2737
rect 580 2731 584 2735
rect 590 2734 594 2738
rect 701 2732 705 2736
rect 719 2733 723 2737
rect 743 2731 747 2735
rect 753 2734 757 2738
rect 857 2732 861 2736
rect 875 2733 879 2737
rect 899 2731 903 2735
rect 909 2734 913 2738
rect 995 2732 999 2736
rect 1013 2733 1017 2737
rect 1037 2731 1041 2735
rect 1047 2734 1051 2738
rect 1138 2732 1142 2736
rect 1156 2733 1160 2737
rect 1180 2731 1184 2735
rect 1190 2734 1194 2738
rect 1301 2732 1305 2736
rect 1319 2733 1323 2737
rect 1343 2731 1347 2735
rect 1353 2734 1357 2738
rect 1457 2732 1461 2736
rect 1475 2733 1479 2737
rect 1499 2731 1503 2735
rect 1509 2734 1513 2738
rect 2360 2707 2364 2711
rect 2435 2707 2439 2711
rect 2445 2707 2449 2711
rect 2461 2713 2465 2717
rect 395 2607 399 2611
rect 413 2608 417 2612
rect 437 2606 441 2610
rect 447 2609 451 2613
rect 538 2607 542 2611
rect 556 2608 560 2612
rect 580 2606 584 2610
rect 590 2609 594 2613
rect 701 2607 705 2611
rect 719 2608 723 2612
rect 743 2606 747 2610
rect 753 2609 757 2613
rect 857 2607 861 2611
rect 875 2608 879 2612
rect 899 2606 903 2610
rect 909 2609 913 2613
rect 995 2607 999 2611
rect 1013 2608 1017 2612
rect 1037 2606 1041 2610
rect 1047 2609 1051 2613
rect 1138 2607 1142 2611
rect 1156 2608 1160 2612
rect 1180 2606 1184 2610
rect 1190 2609 1194 2613
rect 1301 2607 1305 2611
rect 1319 2608 1323 2612
rect 1343 2606 1347 2610
rect 1353 2609 1357 2613
rect 1457 2607 1461 2611
rect 1475 2608 1479 2612
rect 1499 2606 1503 2610
rect 1509 2609 1513 2613
rect 777 2248 781 2252
rect 795 2249 799 2253
rect 819 2247 823 2251
rect 829 2250 833 2254
rect 920 2248 924 2252
rect 938 2249 942 2253
rect 962 2247 966 2251
rect 972 2250 976 2254
rect 1083 2248 1087 2252
rect 1101 2249 1105 2253
rect 1125 2247 1129 2251
rect 1135 2250 1139 2254
rect 1239 2248 1243 2252
rect 1257 2249 1261 2253
rect 1281 2247 1285 2251
rect 1291 2250 1295 2254
rect 2118 2664 2122 2668
rect 2126 2664 2130 2668
rect 2810 2662 2814 2666
rect 2823 2665 2827 2669
rect 2836 2662 2840 2666
rect 2849 2665 2853 2669
rect 2862 2665 2866 2669
rect 2870 2665 2874 2669
rect 2883 2665 2887 2669
rect 2491 2607 2495 2611
rect 2553 2607 2557 2611
rect 2562 2607 2566 2611
rect 2578 2613 2582 2617
rect 2120 2598 2124 2602
rect 2128 2598 2132 2602
rect 2123 2531 2127 2535
rect 2131 2531 2135 2535
rect 2123 2464 2127 2468
rect 2131 2464 2135 2468
rect 2141 2359 2145 2363
rect 2149 2359 2153 2363
rect 2041 2315 2045 2319
rect 2050 2315 2054 2319
rect 2060 2315 2064 2319
rect 2069 2315 2073 2319
rect 2085 2315 2089 2319
rect 2094 2315 2098 2319
rect 2104 2315 2108 2319
rect 2113 2315 2117 2319
rect 2143 2198 2147 2202
rect 2151 2198 2155 2202
rect 2043 2154 2047 2158
rect 2052 2154 2056 2158
rect 2062 2154 2066 2158
rect 2071 2154 2075 2158
rect 2087 2154 2091 2158
rect 2096 2154 2100 2158
rect 2106 2154 2110 2158
rect 2115 2154 2119 2158
rect 2629 2569 2633 2573
rect 2679 2569 2683 2573
rect 2688 2569 2692 2573
rect 2704 2575 2708 2579
rect 2806 2541 2810 2545
rect 2814 2541 2818 2545
rect 2758 2537 2762 2541
rect 2790 2534 2794 2538
rect 2738 2133 2742 2137
rect 2800 2133 2804 2137
rect 2809 2133 2813 2137
rect 2825 2139 2829 2143
rect 2901 2133 2905 2137
rect 2920 2134 2924 2138
rect 2943 2132 2947 2136
rect 2953 2135 2957 2139
rect 2142 2044 2146 2048
rect 2150 2044 2154 2048
rect 2042 2000 2046 2004
rect 2051 2000 2055 2004
rect 2061 2000 2065 2004
rect 2070 2000 2074 2004
rect 2086 2000 2090 2004
rect 2095 2000 2099 2004
rect 2105 2000 2109 2004
rect 2114 2000 2118 2004
rect 2142 1896 2146 1900
rect 2150 1896 2154 1900
rect 2801 1882 2805 1886
rect 2814 1885 2818 1889
rect 2827 1882 2831 1886
rect 2840 1885 2844 1889
rect 2853 1885 2857 1889
rect 2861 1885 2865 1889
rect 2874 1885 2878 1889
rect 2042 1852 2046 1856
rect 2051 1852 2055 1856
rect 2061 1852 2065 1856
rect 2070 1852 2074 1856
rect 2086 1852 2090 1856
rect 2095 1852 2099 1856
rect 2105 1852 2109 1856
rect 2114 1852 2118 1856
rect 2575 1818 2579 1822
rect 2650 1818 2654 1822
rect 2660 1818 2664 1822
rect 2676 1824 2680 1828
rect 2118 1769 2122 1773
rect 2126 1769 2130 1773
rect 2443 1734 2447 1738
rect 2505 1734 2509 1738
rect 2514 1734 2518 1738
rect 2530 1740 2534 1744
rect 2120 1703 2124 1707
rect 2128 1703 2132 1707
rect 2302 1659 2306 1663
rect 2352 1659 2356 1663
rect 2361 1659 2365 1663
rect 2377 1665 2381 1669
rect 2123 1636 2127 1640
rect 2131 1636 2135 1640
rect 2255 1597 2259 1601
rect 2263 1597 2267 1601
rect 2207 1593 2211 1597
rect 2239 1590 2243 1594
rect 2123 1569 2127 1573
rect 2131 1569 2135 1573
<< pdcontact >>
rect 208 3545 212 3549
rect 217 3545 221 3549
rect 234 3545 238 3549
rect 243 3545 247 3549
rect 259 3546 263 3550
rect 269 3545 273 3549
rect 284 3547 288 3551
rect 293 3545 297 3549
rect 385 3546 389 3550
rect 394 3546 398 3550
rect 411 3546 415 3550
rect 420 3546 424 3550
rect 436 3547 440 3551
rect 446 3546 450 3550
rect 461 3548 465 3552
rect 470 3546 474 3550
rect 771 3552 775 3556
rect 780 3552 784 3556
rect 797 3552 801 3556
rect 806 3552 810 3556
rect 822 3553 826 3557
rect 832 3552 836 3556
rect 847 3554 851 3558
rect 856 3552 860 3556
rect 234 3456 238 3460
rect 243 3453 247 3457
rect 252 3456 256 3460
rect 276 3456 280 3460
rect 286 3455 290 3459
rect 948 3553 952 3557
rect 957 3553 961 3557
rect 974 3553 978 3557
rect 983 3553 987 3557
rect 999 3554 1003 3558
rect 1009 3553 1013 3557
rect 1024 3555 1028 3559
rect 1033 3553 1037 3557
rect 1347 3538 1351 3542
rect 1356 3538 1360 3542
rect 1373 3538 1377 3542
rect 1382 3538 1386 3542
rect 1398 3539 1402 3543
rect 1408 3538 1412 3542
rect 1423 3540 1427 3544
rect 1432 3538 1436 3542
rect 550 3469 554 3473
rect 420 3462 424 3466
rect 429 3459 433 3463
rect 438 3462 442 3466
rect 462 3462 466 3466
rect 472 3461 476 3465
rect 573 3466 577 3470
rect 606 3469 610 3473
rect 616 3468 620 3472
rect 797 3463 801 3467
rect 806 3460 810 3464
rect 815 3463 819 3467
rect 839 3463 843 3467
rect 849 3462 853 3466
rect 1113 3476 1117 3480
rect 983 3469 987 3473
rect 992 3466 996 3470
rect 1001 3469 1005 3473
rect 1025 3469 1029 3473
rect 1035 3468 1039 3472
rect 1136 3473 1140 3477
rect 1169 3476 1173 3480
rect 1179 3475 1183 3479
rect 1524 3539 1528 3543
rect 1533 3539 1537 3543
rect 1550 3539 1554 3543
rect 1559 3539 1563 3543
rect 1575 3540 1579 3544
rect 1585 3539 1589 3543
rect 1600 3541 1604 3545
rect 1609 3539 1613 3543
rect 1968 3569 1972 3573
rect 1977 3569 1981 3573
rect 1994 3569 1998 3573
rect 2003 3569 2007 3573
rect 2019 3570 2023 3574
rect 2029 3569 2033 3573
rect 2044 3571 2048 3575
rect 2053 3569 2057 3573
rect 2145 3570 2149 3574
rect 2154 3570 2158 3574
rect 2171 3570 2175 3574
rect 2180 3570 2184 3574
rect 2196 3571 2200 3575
rect 2206 3570 2210 3574
rect 2221 3572 2225 3576
rect 2230 3570 2234 3574
rect 1373 3449 1377 3453
rect 1382 3446 1386 3450
rect 1391 3449 1395 3453
rect 1415 3449 1419 3453
rect 1425 3448 1429 3452
rect 1689 3462 1693 3466
rect 1559 3455 1563 3459
rect 1568 3452 1572 3456
rect 1577 3455 1581 3459
rect 1601 3455 1605 3459
rect 1611 3454 1615 3458
rect 1712 3459 1716 3463
rect 1745 3462 1749 3466
rect 1994 3480 1998 3484
rect 2003 3477 2007 3481
rect 2012 3480 2016 3484
rect 2036 3480 2040 3484
rect 2046 3479 2050 3483
rect 1755 3461 1759 3465
rect 2310 3493 2314 3497
rect 2180 3486 2184 3490
rect 2189 3483 2193 3487
rect 2198 3486 2202 3490
rect 2222 3486 2226 3490
rect 2232 3485 2236 3489
rect 2333 3490 2337 3494
rect 2366 3493 2370 3497
rect 2376 3492 2380 3496
rect 395 3056 399 3060
rect 404 3053 408 3057
rect 413 3056 417 3060
rect 437 3056 441 3060
rect 447 3055 451 3059
rect 538 3056 542 3060
rect 547 3053 551 3057
rect 556 3056 560 3060
rect 580 3056 584 3060
rect 590 3055 594 3059
rect 701 3056 705 3060
rect 710 3053 714 3057
rect 719 3056 723 3060
rect 743 3056 747 3060
rect 753 3055 757 3059
rect 857 3056 861 3060
rect 866 3053 870 3057
rect 875 3056 879 3060
rect 899 3056 903 3060
rect 909 3055 913 3059
rect 995 3056 999 3060
rect 1004 3053 1008 3057
rect 1013 3056 1017 3060
rect 1037 3056 1041 3060
rect 1047 3055 1051 3059
rect 1138 3056 1142 3060
rect 1147 3053 1151 3057
rect 1156 3056 1160 3060
rect 1180 3056 1184 3060
rect 1190 3055 1194 3059
rect 1301 3056 1305 3060
rect 1310 3053 1314 3057
rect 1319 3056 1323 3060
rect 1343 3056 1347 3060
rect 1353 3055 1357 3059
rect 1457 3056 1461 3060
rect 1466 3053 1470 3057
rect 1475 3056 1479 3060
rect 1499 3056 1503 3060
rect 1509 3055 1513 3059
rect 2965 3245 2969 3249
rect 2974 3245 2978 3249
rect 2991 3245 2995 3249
rect 3000 3245 3004 3249
rect 3016 3246 3020 3250
rect 3026 3245 3030 3249
rect 3041 3247 3045 3251
rect 3050 3245 3054 3249
rect 3142 3246 3146 3250
rect 3151 3246 3155 3250
rect 3168 3246 3172 3250
rect 3177 3246 3181 3250
rect 3193 3247 3197 3251
rect 3203 3246 3207 3250
rect 3218 3248 3222 3252
rect 3227 3246 3231 3250
rect 3528 3252 3532 3256
rect 3537 3252 3541 3256
rect 3554 3252 3558 3256
rect 3563 3252 3567 3256
rect 3579 3253 3583 3257
rect 3589 3252 3593 3256
rect 3604 3254 3608 3258
rect 3613 3252 3617 3256
rect 2991 3156 2995 3160
rect 3000 3153 3004 3157
rect 3009 3156 3013 3160
rect 3033 3156 3037 3160
rect 3043 3155 3047 3159
rect 3705 3253 3709 3257
rect 3714 3253 3718 3257
rect 3731 3253 3735 3257
rect 3740 3253 3744 3257
rect 3756 3254 3760 3258
rect 3766 3253 3770 3257
rect 3781 3255 3785 3259
rect 3790 3253 3794 3257
rect 4104 3238 4108 3242
rect 4113 3238 4117 3242
rect 4130 3238 4134 3242
rect 4139 3238 4143 3242
rect 4155 3239 4159 3243
rect 4165 3238 4169 3242
rect 4180 3240 4184 3244
rect 4189 3238 4193 3242
rect 3307 3169 3311 3173
rect 3177 3162 3181 3166
rect 3186 3159 3190 3163
rect 3195 3162 3199 3166
rect 3219 3162 3223 3166
rect 3229 3161 3233 3165
rect 3330 3166 3334 3170
rect 3363 3169 3367 3173
rect 3373 3168 3377 3172
rect 3554 3163 3558 3167
rect 3563 3160 3567 3164
rect 3572 3163 3576 3167
rect 3596 3163 3600 3167
rect 3606 3162 3610 3166
rect 3870 3176 3874 3180
rect 3740 3169 3744 3173
rect 3749 3166 3753 3170
rect 3758 3169 3762 3173
rect 3782 3169 3786 3173
rect 3792 3168 3796 3172
rect 3893 3173 3897 3177
rect 3926 3176 3930 3180
rect 3936 3175 3940 3179
rect 4281 3239 4285 3243
rect 4290 3239 4294 3243
rect 4307 3239 4311 3243
rect 4316 3239 4320 3243
rect 4332 3240 4336 3244
rect 4342 3239 4346 3243
rect 4357 3241 4361 3245
rect 4366 3239 4370 3243
rect 4725 3269 4729 3273
rect 4734 3269 4738 3273
rect 4751 3269 4755 3273
rect 4760 3269 4764 3273
rect 4776 3270 4780 3274
rect 4786 3269 4790 3273
rect 4801 3271 4805 3275
rect 4810 3269 4814 3273
rect 4902 3270 4906 3274
rect 4911 3270 4915 3274
rect 4928 3270 4932 3274
rect 4937 3270 4941 3274
rect 4953 3271 4957 3275
rect 4963 3270 4967 3274
rect 4978 3272 4982 3276
rect 4987 3270 4991 3274
rect 4130 3149 4134 3153
rect 4139 3146 4143 3150
rect 4148 3149 4152 3153
rect 4172 3149 4176 3153
rect 4182 3148 4186 3152
rect 4446 3162 4450 3166
rect 4316 3155 4320 3159
rect 4325 3152 4329 3156
rect 4334 3155 4338 3159
rect 4358 3155 4362 3159
rect 4368 3154 4372 3158
rect 4469 3159 4473 3163
rect 4502 3162 4506 3166
rect 4751 3180 4755 3184
rect 4760 3177 4764 3181
rect 4769 3180 4773 3184
rect 4793 3180 4797 3184
rect 4803 3179 4807 3183
rect 4512 3161 4516 3165
rect 5067 3193 5071 3197
rect 4937 3186 4941 3190
rect 4946 3183 4950 3187
rect 4955 3186 4959 3190
rect 4979 3186 4983 3190
rect 4989 3185 4993 3189
rect 5090 3190 5094 3194
rect 5123 3193 5127 3197
rect 5133 3192 5137 3196
rect 237 2988 241 2992
rect 246 2985 250 2989
rect 255 2988 259 2992
rect 279 2988 283 2992
rect 289 2987 293 2991
rect 189 2934 193 2938
rect 197 2934 201 2938
rect 100 2904 104 2908
rect 109 2901 113 2905
rect 118 2904 122 2908
rect 142 2904 146 2908
rect 152 2903 156 2907
rect 236 2907 240 2911
rect 245 2904 249 2908
rect 254 2907 258 2911
rect 278 2907 282 2911
rect 288 2906 292 2910
rect 189 2851 193 2855
rect 197 2851 201 2855
rect 395 2914 399 2918
rect 404 2911 408 2915
rect 413 2914 417 2918
rect 437 2914 441 2918
rect 447 2913 451 2917
rect 538 2914 542 2918
rect 547 2911 551 2915
rect 556 2914 560 2918
rect 580 2914 584 2918
rect 590 2913 594 2917
rect 701 2914 705 2918
rect 710 2911 714 2915
rect 719 2914 723 2918
rect 743 2914 747 2918
rect 753 2913 757 2917
rect 857 2914 861 2918
rect 866 2911 870 2915
rect 875 2914 879 2918
rect 899 2914 903 2918
rect 909 2913 913 2917
rect 995 2914 999 2918
rect 1004 2911 1008 2915
rect 1013 2914 1017 2918
rect 1037 2914 1041 2918
rect 1047 2913 1051 2917
rect 1138 2914 1142 2918
rect 1147 2911 1151 2915
rect 1156 2914 1160 2918
rect 1180 2914 1184 2918
rect 1190 2913 1194 2917
rect 1301 2914 1305 2918
rect 1310 2911 1314 2915
rect 1319 2914 1323 2918
rect 1343 2914 1347 2918
rect 1353 2913 1357 2917
rect 1457 2914 1461 2918
rect 1466 2911 1470 2915
rect 1475 2914 1479 2918
rect 1499 2914 1503 2918
rect 1509 2913 1513 2917
rect 1692 2935 1696 2939
rect 1701 2935 1705 2939
rect 1718 2935 1722 2939
rect 1727 2935 1731 2939
rect 1743 2936 1747 2940
rect 1753 2935 1757 2939
rect 1768 2937 1772 2941
rect 1777 2935 1781 2939
rect 1887 2936 1891 2940
rect 1896 2936 1900 2940
rect 1913 2936 1917 2940
rect 1922 2936 1926 2940
rect 1938 2937 1942 2941
rect 1948 2936 1952 2940
rect 1963 2938 1967 2942
rect 1972 2936 1976 2940
rect 2100 2935 2104 2939
rect 2109 2935 2113 2939
rect 2126 2935 2130 2939
rect 2135 2935 2139 2939
rect 2151 2936 2155 2940
rect 2161 2935 2165 2939
rect 2176 2937 2180 2941
rect 2185 2935 2189 2939
rect 2301 2936 2305 2940
rect 2310 2936 2314 2940
rect 2327 2936 2331 2940
rect 2336 2936 2340 2940
rect 2352 2937 2356 2941
rect 2362 2936 2366 2940
rect 2377 2938 2381 2942
rect 2386 2936 2390 2940
rect 240 2816 244 2820
rect 249 2813 253 2817
rect 258 2816 262 2820
rect 282 2816 286 2820
rect 292 2815 296 2819
rect 395 2765 399 2769
rect 404 2762 408 2766
rect 413 2765 417 2769
rect 437 2765 441 2769
rect 447 2764 451 2768
rect 538 2765 542 2769
rect 547 2762 551 2766
rect 556 2765 560 2769
rect 580 2765 584 2769
rect 590 2764 594 2768
rect 701 2765 705 2769
rect 710 2762 714 2766
rect 719 2765 723 2769
rect 743 2765 747 2769
rect 753 2764 757 2768
rect 857 2765 861 2769
rect 866 2762 870 2766
rect 875 2765 879 2769
rect 899 2765 903 2769
rect 909 2764 913 2768
rect 995 2765 999 2769
rect 1004 2762 1008 2766
rect 1013 2765 1017 2769
rect 1037 2765 1041 2769
rect 1047 2764 1051 2768
rect 1138 2765 1142 2769
rect 1147 2762 1151 2766
rect 1156 2765 1160 2769
rect 1180 2765 1184 2769
rect 1190 2764 1194 2768
rect 1301 2765 1305 2769
rect 1310 2762 1314 2766
rect 1319 2765 1323 2769
rect 1343 2765 1347 2769
rect 1353 2764 1357 2768
rect 1457 2765 1461 2769
rect 1466 2762 1470 2766
rect 1475 2765 1479 2769
rect 1499 2765 1503 2769
rect 1509 2764 1513 2768
rect 2360 2742 2364 2746
rect 2373 2742 2377 2746
rect 2390 2742 2394 2746
rect 2405 2742 2409 2746
rect 2420 2742 2424 2746
rect 2435 2742 2439 2746
rect 2445 2742 2449 2746
rect 2461 2742 2465 2746
rect 2118 2688 2122 2692
rect 2126 2688 2130 2692
rect 395 2640 399 2644
rect 404 2637 408 2641
rect 413 2640 417 2644
rect 437 2640 441 2644
rect 447 2639 451 2643
rect 538 2640 542 2644
rect 547 2637 551 2641
rect 556 2640 560 2644
rect 580 2640 584 2644
rect 590 2639 594 2643
rect 701 2640 705 2644
rect 710 2637 714 2641
rect 719 2640 723 2644
rect 743 2640 747 2644
rect 753 2639 757 2643
rect 857 2640 861 2644
rect 866 2637 870 2641
rect 875 2640 879 2644
rect 899 2640 903 2644
rect 909 2639 913 2643
rect 995 2640 999 2644
rect 1004 2637 1008 2641
rect 1013 2640 1017 2644
rect 1037 2640 1041 2644
rect 1047 2639 1051 2643
rect 1138 2640 1142 2644
rect 1147 2637 1151 2641
rect 1156 2640 1160 2644
rect 1180 2640 1184 2644
rect 1190 2639 1194 2643
rect 1301 2640 1305 2644
rect 1310 2637 1314 2641
rect 1319 2640 1323 2644
rect 1343 2640 1347 2644
rect 1353 2639 1357 2643
rect 1457 2640 1461 2644
rect 1466 2637 1470 2641
rect 1475 2640 1479 2644
rect 1499 2640 1503 2644
rect 1509 2639 1513 2643
rect 777 2281 781 2285
rect 786 2278 790 2282
rect 795 2281 799 2285
rect 819 2281 823 2285
rect 829 2280 833 2284
rect 920 2281 924 2285
rect 929 2278 933 2282
rect 938 2281 942 2285
rect 962 2281 966 2285
rect 972 2280 976 2284
rect 1083 2281 1087 2285
rect 1092 2278 1096 2282
rect 1101 2281 1105 2285
rect 1125 2281 1129 2285
rect 1135 2280 1139 2284
rect 1239 2281 1243 2285
rect 1248 2278 1252 2282
rect 1257 2281 1261 2285
rect 1281 2281 1285 2285
rect 1291 2280 1295 2284
rect 2491 2642 2495 2646
rect 2506 2642 2511 2646
rect 2524 2642 2528 2646
rect 2539 2642 2543 2646
rect 2553 2642 2557 2646
rect 2562 2642 2566 2646
rect 2578 2642 2582 2646
rect 2810 2692 2814 2696
rect 2862 2692 2866 2696
rect 2870 2692 2874 2696
rect 2883 2692 2887 2696
rect 2120 2622 2124 2626
rect 2128 2622 2132 2626
rect 2123 2555 2127 2559
rect 2131 2555 2135 2559
rect 2123 2488 2127 2492
rect 2131 2488 2135 2492
rect 2141 2383 2145 2387
rect 2149 2383 2153 2387
rect 2041 2346 2045 2350
rect 2050 2346 2054 2350
rect 2060 2346 2064 2350
rect 2069 2346 2073 2350
rect 2085 2346 2089 2350
rect 2094 2346 2098 2350
rect 2104 2346 2108 2350
rect 2113 2346 2117 2350
rect 2143 2222 2147 2226
rect 2151 2222 2155 2226
rect 2043 2185 2047 2189
rect 2052 2185 2056 2189
rect 2062 2185 2066 2189
rect 2071 2185 2075 2189
rect 2087 2185 2091 2189
rect 2096 2185 2100 2189
rect 2106 2185 2110 2189
rect 2115 2185 2119 2189
rect 2629 2604 2633 2608
rect 2644 2604 2649 2608
rect 2662 2604 2666 2608
rect 2679 2604 2683 2608
rect 2688 2604 2692 2608
rect 2704 2604 2708 2608
rect 2758 2564 2762 2568
rect 2769 2565 2773 2569
rect 2779 2564 2783 2568
rect 2790 2565 2794 2569
rect 2806 2565 2810 2569
rect 2814 2565 2818 2569
rect 2738 2168 2742 2172
rect 2753 2168 2758 2172
rect 2771 2168 2775 2172
rect 2786 2168 2790 2172
rect 2800 2168 2804 2172
rect 2809 2168 2813 2172
rect 2825 2168 2829 2172
rect 2901 2166 2905 2170
rect 2912 2163 2916 2167
rect 2921 2166 2925 2170
rect 2943 2166 2947 2170
rect 2953 2165 2957 2169
rect 2142 2068 2146 2072
rect 2150 2068 2154 2072
rect 2042 2031 2046 2035
rect 2051 2031 2055 2035
rect 2061 2031 2065 2035
rect 2070 2031 2074 2035
rect 2086 2031 2090 2035
rect 2095 2031 2099 2035
rect 2105 2031 2109 2035
rect 2114 2031 2118 2035
rect 2142 1920 2146 1924
rect 2150 1920 2154 1924
rect 2801 1912 2805 1916
rect 2853 1912 2857 1916
rect 2861 1912 2865 1916
rect 2874 1912 2878 1916
rect 2042 1883 2046 1887
rect 2051 1883 2055 1887
rect 2061 1883 2065 1887
rect 2070 1883 2074 1887
rect 2086 1883 2090 1887
rect 2095 1883 2099 1887
rect 2105 1883 2109 1887
rect 2114 1883 2118 1887
rect 2575 1853 2579 1857
rect 2588 1853 2592 1857
rect 2605 1853 2609 1857
rect 2620 1853 2624 1857
rect 2635 1853 2639 1857
rect 2650 1853 2654 1857
rect 2660 1853 2664 1857
rect 2676 1853 2680 1857
rect 2118 1793 2122 1797
rect 2126 1793 2130 1797
rect 2443 1769 2447 1773
rect 2458 1769 2463 1773
rect 2476 1769 2480 1773
rect 2491 1769 2495 1773
rect 2505 1769 2509 1773
rect 2514 1769 2518 1773
rect 2530 1769 2534 1773
rect 2120 1727 2124 1731
rect 2128 1727 2132 1731
rect 2302 1694 2306 1698
rect 2317 1694 2322 1698
rect 2335 1694 2339 1698
rect 2352 1694 2356 1698
rect 2361 1694 2365 1698
rect 2377 1694 2381 1698
rect 2123 1660 2127 1664
rect 2131 1660 2135 1664
rect 2207 1620 2211 1624
rect 2218 1621 2222 1625
rect 2228 1620 2232 1624
rect 2239 1621 2243 1625
rect 2255 1621 2259 1625
rect 2263 1621 2267 1625
rect 2123 1593 2127 1597
rect 2131 1593 2135 1597
<< polysilicon >>
rect 25 3731 208 3732
rect 24 3723 208 3731
rect 24 3690 30 3723
rect 794 3732 801 3733
rect 220 3723 2466 3732
rect 24 3074 31 3690
rect 794 3649 801 3723
rect 1335 3626 1341 3723
rect 1986 3657 1991 3723
rect 1335 3617 1341 3618
rect 1993 3605 2095 3608
rect 1018 3594 1033 3597
rect 455 3587 475 3590
rect 233 3581 335 3584
rect 233 3571 236 3581
rect 264 3571 322 3574
rect 198 3560 241 3562
rect 198 3504 200 3560
rect 213 3550 215 3555
rect 239 3550 241 3560
rect 264 3550 266 3571
rect 290 3550 292 3554
rect 213 3536 215 3545
rect 239 3542 241 3545
rect 213 3534 241 3536
rect 213 3519 215 3522
rect 239 3519 241 3534
rect 264 3533 266 3545
rect 264 3519 266 3529
rect 290 3519 292 3545
rect 300 3531 306 3533
rect 213 3504 215 3514
rect 198 3502 215 3504
rect 213 3497 215 3502
rect 239 3503 241 3514
rect 264 3511 266 3514
rect 239 3501 245 3503
rect 290 3503 292 3514
rect 249 3501 292 3503
rect 304 3497 306 3531
rect 213 3495 306 3497
rect 319 3472 322 3571
rect 406 3571 409 3585
rect 375 3561 418 3563
rect 375 3505 377 3561
rect 390 3551 392 3556
rect 416 3551 418 3561
rect 441 3551 443 3554
rect 390 3537 392 3546
rect 416 3543 418 3546
rect 441 3537 443 3546
rect 455 3537 458 3587
rect 482 3587 501 3590
rect 467 3551 469 3555
rect 390 3535 418 3537
rect 390 3520 392 3523
rect 416 3520 418 3535
rect 441 3535 458 3537
rect 441 3534 443 3535
rect 441 3520 443 3530
rect 467 3520 469 3546
rect 477 3532 483 3534
rect 390 3505 392 3515
rect 375 3503 392 3505
rect 390 3498 392 3503
rect 416 3504 418 3515
rect 441 3512 443 3515
rect 416 3502 438 3504
rect 467 3504 469 3515
rect 442 3502 469 3504
rect 481 3498 483 3532
rect 390 3496 483 3498
rect 497 3486 501 3587
rect 796 3588 898 3591
rect 796 3578 799 3588
rect 827 3578 885 3581
rect 761 3567 804 3569
rect 761 3511 763 3567
rect 776 3557 778 3562
rect 802 3557 804 3567
rect 827 3557 829 3578
rect 853 3557 855 3561
rect 776 3543 778 3552
rect 802 3549 804 3552
rect 776 3541 804 3543
rect 776 3526 778 3529
rect 802 3526 804 3541
rect 827 3540 829 3552
rect 827 3526 829 3536
rect 853 3526 855 3552
rect 863 3538 869 3540
rect 776 3511 778 3521
rect 761 3509 778 3511
rect 776 3504 778 3509
rect 802 3510 804 3521
rect 827 3518 829 3521
rect 802 3508 808 3510
rect 853 3510 855 3521
rect 812 3508 855 3510
rect 867 3504 869 3538
rect 776 3502 869 3504
rect 218 3469 322 3472
rect 397 3483 501 3486
rect 218 3464 221 3469
rect 218 3443 221 3458
rect 239 3459 241 3462
rect 248 3459 250 3462
rect 239 3443 241 3454
rect 281 3459 283 3462
rect 218 3440 241 3443
rect 239 3428 241 3440
rect 248 3435 250 3454
rect 281 3443 283 3454
rect 397 3449 400 3483
rect 882 3479 885 3578
rect 969 3578 972 3588
rect 938 3568 981 3570
rect 938 3512 940 3568
rect 953 3558 955 3563
rect 979 3558 981 3568
rect 1004 3558 1006 3561
rect 953 3544 955 3553
rect 979 3550 981 3553
rect 1004 3544 1006 3553
rect 1018 3544 1021 3594
rect 1039 3594 1064 3597
rect 1993 3595 1996 3605
rect 1030 3558 1032 3562
rect 953 3542 981 3544
rect 953 3527 955 3530
rect 979 3527 981 3542
rect 1004 3542 1021 3544
rect 1004 3541 1006 3542
rect 1004 3527 1006 3537
rect 1030 3527 1032 3553
rect 1040 3539 1046 3541
rect 953 3512 955 3522
rect 938 3510 955 3512
rect 953 3505 955 3510
rect 979 3511 981 3522
rect 1004 3519 1006 3522
rect 979 3509 1001 3511
rect 1030 3511 1032 3522
rect 1005 3509 1032 3511
rect 1044 3505 1046 3539
rect 953 3503 1046 3505
rect 1060 3493 1064 3594
rect 2024 3595 2082 3598
rect 1594 3580 1619 3583
rect 1372 3574 1474 3577
rect 1372 3564 1375 3574
rect 1403 3564 1461 3567
rect 1337 3553 1380 3555
rect 1337 3497 1339 3553
rect 1352 3543 1354 3548
rect 1378 3543 1380 3553
rect 1403 3543 1405 3564
rect 1429 3543 1431 3547
rect 1352 3529 1354 3538
rect 1378 3535 1380 3538
rect 1352 3527 1380 3529
rect 1352 3512 1354 3515
rect 1378 3512 1380 3527
rect 1403 3526 1405 3538
rect 1403 3512 1405 3522
rect 1429 3512 1431 3538
rect 1439 3524 1445 3526
rect 1352 3497 1354 3507
rect 1337 3495 1354 3497
rect 779 3476 885 3479
rect 960 3490 1064 3493
rect 1352 3490 1354 3495
rect 1378 3496 1380 3507
rect 1403 3504 1405 3507
rect 1378 3494 1384 3496
rect 1429 3496 1431 3507
rect 1388 3494 1431 3496
rect 1443 3490 1445 3524
rect 555 3472 557 3475
rect 565 3472 567 3475
rect 425 3465 427 3468
rect 434 3465 436 3468
rect 425 3449 427 3460
rect 467 3465 469 3468
rect 397 3446 427 3449
rect 282 3439 283 3443
rect 249 3431 250 3435
rect 248 3428 250 3431
rect 281 3428 283 3439
rect 425 3434 427 3446
rect 434 3441 436 3460
rect 467 3449 469 3460
rect 435 3437 436 3441
rect 434 3434 436 3437
rect 467 3434 469 3445
rect 239 3420 241 3423
rect 248 3420 250 3423
rect 425 3426 427 3429
rect 434 3426 436 3429
rect 467 3426 469 3429
rect 281 3420 283 3423
rect 535 3406 539 3452
rect 555 3447 557 3467
rect 565 3456 567 3467
rect 611 3472 613 3475
rect 779 3467 782 3476
rect 555 3433 557 3443
rect 565 3433 567 3452
rect 611 3448 613 3467
rect 612 3444 613 3448
rect 779 3450 782 3462
rect 802 3466 804 3469
rect 811 3466 813 3469
rect 802 3450 804 3461
rect 844 3466 846 3469
rect 779 3447 804 3450
rect 611 3433 613 3444
rect 802 3435 804 3447
rect 811 3442 813 3461
rect 844 3450 846 3461
rect 960 3456 963 3490
rect 1352 3488 1445 3490
rect 1118 3479 1120 3482
rect 1128 3479 1130 3482
rect 988 3472 990 3475
rect 997 3472 999 3475
rect 988 3456 990 3467
rect 1030 3472 1032 3475
rect 960 3453 990 3456
rect 845 3446 846 3450
rect 812 3438 813 3442
rect 811 3435 813 3438
rect 844 3435 846 3446
rect 988 3441 990 3453
rect 997 3448 999 3467
rect 1030 3456 1032 3467
rect 998 3444 999 3448
rect 997 3441 999 3444
rect 1030 3441 1032 3452
rect 555 3425 557 3428
rect 565 3425 567 3428
rect 611 3425 613 3428
rect 802 3427 804 3430
rect 811 3427 813 3430
rect 988 3433 990 3436
rect 997 3433 999 3436
rect 1030 3433 1032 3436
rect 844 3427 846 3430
rect 1098 3413 1102 3459
rect 1118 3454 1120 3474
rect 1128 3463 1130 3474
rect 1174 3479 1176 3482
rect 1118 3440 1120 3450
rect 1128 3440 1130 3459
rect 1174 3455 1176 3474
rect 1458 3465 1461 3564
rect 1545 3564 1548 3574
rect 1514 3554 1557 3556
rect 1514 3498 1516 3554
rect 1529 3544 1531 3549
rect 1555 3544 1557 3554
rect 1580 3544 1582 3547
rect 1529 3530 1531 3539
rect 1555 3536 1557 3539
rect 1580 3530 1582 3539
rect 1594 3530 1597 3580
rect 1958 3584 2001 3586
rect 1627 3580 1640 3583
rect 1606 3544 1608 3548
rect 1529 3528 1557 3530
rect 1529 3513 1531 3516
rect 1555 3513 1557 3528
rect 1580 3528 1597 3530
rect 1580 3527 1582 3528
rect 1580 3513 1582 3523
rect 1606 3513 1608 3539
rect 1616 3525 1622 3527
rect 1529 3498 1531 3508
rect 1514 3496 1531 3498
rect 1529 3491 1531 3496
rect 1555 3497 1557 3508
rect 1580 3505 1582 3508
rect 1555 3495 1577 3497
rect 1606 3497 1608 3508
rect 1581 3495 1608 3497
rect 1620 3491 1622 3525
rect 1529 3489 1622 3491
rect 1636 3479 1640 3580
rect 1958 3528 1960 3584
rect 1973 3574 1975 3579
rect 1999 3574 2001 3584
rect 2024 3574 2026 3595
rect 2050 3574 2052 3578
rect 1973 3560 1975 3569
rect 1999 3566 2001 3569
rect 1973 3558 2001 3560
rect 1973 3543 1975 3546
rect 1999 3543 2001 3558
rect 2024 3557 2026 3569
rect 2024 3543 2026 3553
rect 2050 3543 2052 3569
rect 2060 3555 2066 3557
rect 1973 3528 1975 3538
rect 1958 3526 1975 3528
rect 1973 3521 1975 3526
rect 1999 3527 2001 3538
rect 2024 3535 2026 3538
rect 1999 3525 2005 3527
rect 2050 3527 2052 3538
rect 2009 3525 2052 3527
rect 2064 3521 2066 3555
rect 1973 3519 2066 3521
rect 2079 3496 2082 3595
rect 2166 3595 2169 3613
rect 2215 3611 2261 3614
rect 2135 3585 2178 3587
rect 2135 3529 2137 3585
rect 2150 3575 2152 3580
rect 2176 3575 2178 3585
rect 2201 3575 2203 3578
rect 2150 3561 2152 3570
rect 2176 3567 2178 3570
rect 2201 3561 2203 3570
rect 2215 3561 2218 3611
rect 2227 3575 2229 3579
rect 2150 3559 2178 3561
rect 2150 3544 2152 3547
rect 2176 3544 2178 3559
rect 2201 3559 2218 3561
rect 2201 3558 2203 3559
rect 2201 3544 2203 3554
rect 2227 3544 2229 3570
rect 2257 3564 2261 3611
rect 2237 3556 2243 3558
rect 2150 3529 2152 3539
rect 2135 3527 2152 3529
rect 2150 3522 2152 3527
rect 2176 3528 2178 3539
rect 2201 3536 2203 3539
rect 2176 3526 2198 3528
rect 2227 3528 2229 3539
rect 2202 3526 2229 3528
rect 2241 3522 2243 3556
rect 2150 3520 2243 3522
rect 2257 3510 2261 3557
rect 1968 3493 2082 3496
rect 2157 3507 2261 3510
rect 1175 3451 1176 3455
rect 1174 3440 1176 3451
rect 1353 3462 1461 3465
rect 1536 3476 1640 3479
rect 1353 3452 1356 3462
rect 1378 3452 1380 3455
rect 1387 3452 1389 3455
rect 1118 3432 1120 3435
rect 1128 3432 1130 3435
rect 1353 3436 1356 3446
rect 1378 3436 1380 3447
rect 1420 3452 1422 3455
rect 1174 3432 1176 3435
rect 1353 3433 1380 3436
rect 1378 3421 1380 3433
rect 1387 3428 1389 3447
rect 1420 3436 1422 3447
rect 1536 3442 1539 3476
rect 1694 3465 1696 3468
rect 1704 3465 1706 3468
rect 1564 3458 1566 3461
rect 1573 3458 1575 3461
rect 1564 3442 1566 3453
rect 1606 3458 1608 3461
rect 1536 3439 1566 3442
rect 1421 3432 1422 3436
rect 1388 3424 1389 3428
rect 1387 3421 1389 3424
rect 1420 3421 1422 3432
rect 1564 3427 1566 3439
rect 1573 3434 1575 3453
rect 1606 3442 1608 3453
rect 1574 3430 1575 3434
rect 1573 3427 1575 3430
rect 1606 3427 1608 3438
rect 1378 3413 1380 3416
rect 1387 3413 1389 3416
rect 1564 3419 1566 3422
rect 1573 3419 1575 3422
rect 1606 3419 1608 3422
rect 1420 3413 1422 3416
rect 884 3409 1102 3413
rect 321 3402 539 3406
rect 1674 3399 1678 3445
rect 1694 3440 1696 3460
rect 1704 3449 1706 3460
rect 1750 3465 1752 3468
rect 1968 3467 1971 3486
rect 1999 3483 2001 3486
rect 2008 3483 2010 3486
rect 1999 3467 2001 3478
rect 2041 3483 2043 3486
rect 1968 3464 2001 3467
rect 1694 3426 1696 3436
rect 1704 3426 1706 3445
rect 1750 3441 1752 3460
rect 1999 3452 2001 3464
rect 2008 3459 2010 3478
rect 2041 3467 2043 3478
rect 2157 3473 2160 3507
rect 2315 3496 2317 3499
rect 2325 3496 2327 3499
rect 2185 3489 2187 3492
rect 2194 3489 2196 3492
rect 2185 3473 2187 3484
rect 2227 3489 2229 3492
rect 2157 3470 2187 3473
rect 2042 3463 2043 3467
rect 2009 3455 2010 3459
rect 2008 3452 2010 3455
rect 2041 3452 2043 3463
rect 2185 3458 2187 3470
rect 2194 3465 2196 3484
rect 2227 3473 2229 3484
rect 2195 3461 2196 3465
rect 2194 3458 2196 3461
rect 2227 3458 2229 3469
rect 1999 3444 2001 3447
rect 2008 3444 2010 3447
rect 2185 3450 2187 3453
rect 2194 3450 2196 3453
rect 2227 3450 2229 3453
rect 2041 3444 2043 3447
rect 1751 3437 1752 3441
rect 1750 3426 1752 3437
rect 1694 3418 1696 3421
rect 1704 3418 1706 3421
rect 2295 3430 2299 3476
rect 2315 3471 2317 3491
rect 2325 3480 2327 3491
rect 2371 3496 2373 3499
rect 2315 3457 2317 3467
rect 2325 3457 2327 3476
rect 2371 3472 2373 3491
rect 2372 3468 2373 3472
rect 2371 3457 2373 3468
rect 2315 3449 2317 3452
rect 2325 3449 2327 3452
rect 2371 3449 2373 3452
rect 2782 3431 2965 3432
rect 2081 3426 2299 3430
rect 2781 3423 2965 3431
rect 1750 3418 1752 3421
rect 1460 3395 1678 3399
rect 2781 3390 2787 3423
rect 3551 3432 3558 3433
rect 2977 3423 5223 3432
rect 196 3345 415 3352
rect 423 3345 902 3352
rect 2086 3352 2093 3367
rect 910 3345 1556 3352
rect 1564 3346 2093 3352
rect 1564 3345 2092 3346
rect 24 3071 1491 3074
rect 24 3068 310 3071
rect 179 3001 271 3004
rect 58 2949 169 2952
rect 58 2864 62 2949
rect 179 2945 183 3001
rect 268 2999 271 3001
rect 305 3000 309 3068
rect 426 3067 429 3071
rect 569 3067 572 3071
rect 731 3070 735 3071
rect 886 3070 891 3071
rect 732 3067 735 3070
rect 888 3067 891 3070
rect 1026 3067 1029 3071
rect 1169 3067 1172 3071
rect 1331 3070 1335 3071
rect 1332 3067 1335 3070
rect 1488 3067 1491 3071
rect 400 3059 402 3062
rect 409 3059 411 3062
rect 400 3044 402 3054
rect 442 3059 444 3062
rect 543 3059 545 3062
rect 552 3059 554 3062
rect 401 3040 402 3044
rect 400 3028 402 3040
rect 409 3035 411 3054
rect 442 3043 444 3054
rect 543 3044 545 3054
rect 585 3059 587 3062
rect 706 3059 708 3062
rect 715 3059 717 3062
rect 443 3039 444 3043
rect 544 3040 545 3044
rect 410 3031 411 3035
rect 409 3028 411 3031
rect 442 3028 444 3039
rect 400 3020 402 3023
rect 409 3020 411 3023
rect 543 3028 545 3040
rect 552 3035 554 3054
rect 585 3043 587 3054
rect 706 3044 708 3054
rect 748 3059 750 3062
rect 862 3059 864 3062
rect 871 3059 873 3062
rect 586 3039 587 3043
rect 707 3040 708 3044
rect 553 3031 554 3035
rect 552 3028 554 3031
rect 585 3028 587 3039
rect 442 3020 444 3023
rect 543 3020 545 3023
rect 552 3020 554 3023
rect 706 3028 708 3040
rect 715 3035 717 3054
rect 748 3043 750 3054
rect 862 3044 864 3054
rect 904 3059 906 3062
rect 1000 3059 1002 3062
rect 1009 3059 1011 3062
rect 749 3039 750 3043
rect 863 3040 864 3044
rect 716 3031 717 3035
rect 715 3028 717 3031
rect 748 3028 750 3039
rect 585 3020 587 3023
rect 706 3020 708 3023
rect 715 3020 717 3023
rect 862 3028 864 3040
rect 871 3035 873 3054
rect 904 3043 906 3054
rect 1000 3044 1002 3054
rect 1042 3059 1044 3062
rect 1143 3059 1145 3062
rect 1152 3059 1154 3062
rect 905 3039 906 3043
rect 1001 3040 1002 3044
rect 872 3031 873 3035
rect 871 3028 873 3031
rect 904 3028 906 3039
rect 748 3020 750 3023
rect 862 3020 864 3023
rect 871 3020 873 3023
rect 1000 3028 1002 3040
rect 1009 3035 1011 3054
rect 1042 3043 1044 3054
rect 1143 3044 1145 3054
rect 1185 3059 1187 3062
rect 1306 3059 1308 3062
rect 1315 3059 1317 3062
rect 1043 3039 1044 3043
rect 1144 3040 1145 3044
rect 1010 3031 1011 3035
rect 1009 3028 1011 3031
rect 1042 3028 1044 3039
rect 904 3020 906 3023
rect 1000 3020 1002 3023
rect 1009 3020 1011 3023
rect 1143 3028 1145 3040
rect 1152 3035 1154 3054
rect 1185 3043 1187 3054
rect 1306 3044 1308 3054
rect 1348 3059 1350 3062
rect 1462 3059 1464 3062
rect 1471 3059 1473 3062
rect 1186 3039 1187 3043
rect 1307 3040 1308 3044
rect 1153 3031 1154 3035
rect 1152 3028 1154 3031
rect 1185 3028 1187 3039
rect 1042 3020 1044 3023
rect 1143 3020 1145 3023
rect 1152 3020 1154 3023
rect 1306 3028 1308 3040
rect 1315 3035 1317 3054
rect 1348 3043 1350 3054
rect 1462 3044 1464 3054
rect 1504 3059 1506 3062
rect 1349 3039 1350 3043
rect 1463 3040 1464 3044
rect 1316 3031 1317 3035
rect 1315 3028 1317 3031
rect 1348 3028 1350 3039
rect 1185 3020 1187 3023
rect 1306 3020 1308 3023
rect 1315 3020 1317 3023
rect 1462 3028 1464 3040
rect 1471 3035 1473 3054
rect 1504 3043 1506 3054
rect 1505 3039 1506 3043
rect 1472 3031 1473 3035
rect 1471 3028 1473 3031
rect 1504 3028 1506 3039
rect 1348 3020 1350 3023
rect 1462 3020 1464 3023
rect 1471 3020 1473 3023
rect 1504 3020 1506 3023
rect 1539 3008 1541 3013
rect 2085 3013 2092 3345
rect 2781 3029 2788 3390
rect 3551 3349 3558 3423
rect 4092 3326 4098 3423
rect 4743 3357 4748 3423
rect 4092 3317 4098 3318
rect 5014 3314 5020 3388
rect 4750 3305 4852 3308
rect 3775 3294 3790 3297
rect 3212 3287 3232 3290
rect 2990 3281 3092 3284
rect 2990 3271 2993 3281
rect 3021 3271 3079 3274
rect 2955 3260 2998 3262
rect 2955 3204 2957 3260
rect 2970 3250 2972 3255
rect 2996 3250 2998 3260
rect 3021 3250 3023 3271
rect 3047 3250 3049 3254
rect 2970 3236 2972 3245
rect 2996 3242 2998 3245
rect 2970 3234 2998 3236
rect 2970 3219 2972 3222
rect 2996 3219 2998 3234
rect 3021 3233 3023 3245
rect 3021 3219 3023 3229
rect 3047 3219 3049 3245
rect 3057 3231 3063 3233
rect 2970 3204 2972 3214
rect 2955 3202 2972 3204
rect 2970 3197 2972 3202
rect 2996 3203 2998 3214
rect 3021 3211 3023 3214
rect 2996 3201 3002 3203
rect 3047 3203 3049 3214
rect 3006 3201 3049 3203
rect 3061 3197 3063 3231
rect 2970 3195 3063 3197
rect 3076 3172 3079 3271
rect 3163 3271 3166 3285
rect 3132 3261 3175 3263
rect 3132 3205 3134 3261
rect 3147 3251 3149 3256
rect 3173 3251 3175 3261
rect 3198 3251 3200 3254
rect 3147 3237 3149 3246
rect 3173 3243 3175 3246
rect 3198 3237 3200 3246
rect 3212 3237 3215 3287
rect 3239 3287 3258 3290
rect 3224 3251 3226 3255
rect 3147 3235 3175 3237
rect 3147 3220 3149 3223
rect 3173 3220 3175 3235
rect 3198 3235 3215 3237
rect 3198 3234 3200 3235
rect 3198 3220 3200 3230
rect 3224 3220 3226 3246
rect 3234 3232 3240 3234
rect 3147 3205 3149 3215
rect 3132 3203 3149 3205
rect 3147 3198 3149 3203
rect 3173 3204 3175 3215
rect 3198 3212 3200 3215
rect 3173 3202 3195 3204
rect 3224 3204 3226 3215
rect 3199 3202 3226 3204
rect 3238 3198 3240 3232
rect 3147 3196 3240 3198
rect 3254 3186 3258 3287
rect 3553 3288 3655 3291
rect 3553 3278 3556 3288
rect 3584 3278 3642 3281
rect 3518 3267 3561 3269
rect 3518 3211 3520 3267
rect 3533 3257 3535 3262
rect 3559 3257 3561 3267
rect 3584 3257 3586 3278
rect 3610 3257 3612 3261
rect 3533 3243 3535 3252
rect 3559 3249 3561 3252
rect 3533 3241 3561 3243
rect 3533 3226 3535 3229
rect 3559 3226 3561 3241
rect 3584 3240 3586 3252
rect 3584 3226 3586 3236
rect 3610 3226 3612 3252
rect 3620 3238 3626 3240
rect 3533 3211 3535 3221
rect 3518 3209 3535 3211
rect 3533 3204 3535 3209
rect 3559 3210 3561 3221
rect 3584 3218 3586 3221
rect 3559 3208 3565 3210
rect 3610 3210 3612 3221
rect 3569 3208 3612 3210
rect 3624 3204 3626 3238
rect 3533 3202 3626 3204
rect 2975 3169 3079 3172
rect 3154 3183 3258 3186
rect 2975 3164 2978 3169
rect 2975 3143 2978 3158
rect 2996 3159 2998 3162
rect 3005 3159 3007 3162
rect 2996 3143 2998 3154
rect 3038 3159 3040 3162
rect 2975 3140 2998 3143
rect 2996 3128 2998 3140
rect 3005 3135 3007 3154
rect 3038 3143 3040 3154
rect 3154 3149 3157 3183
rect 3639 3179 3642 3278
rect 3726 3278 3729 3288
rect 3695 3268 3738 3270
rect 3695 3212 3697 3268
rect 3710 3258 3712 3263
rect 3736 3258 3738 3268
rect 3761 3258 3763 3261
rect 3710 3244 3712 3253
rect 3736 3250 3738 3253
rect 3761 3244 3763 3253
rect 3775 3244 3778 3294
rect 3796 3294 3821 3297
rect 4750 3295 4753 3305
rect 3787 3258 3789 3262
rect 3710 3242 3738 3244
rect 3710 3227 3712 3230
rect 3736 3227 3738 3242
rect 3761 3242 3778 3244
rect 3761 3241 3763 3242
rect 3761 3227 3763 3237
rect 3787 3227 3789 3253
rect 3797 3239 3803 3241
rect 3710 3212 3712 3222
rect 3695 3210 3712 3212
rect 3710 3205 3712 3210
rect 3736 3211 3738 3222
rect 3761 3219 3763 3222
rect 3736 3209 3758 3211
rect 3787 3211 3789 3222
rect 3762 3209 3789 3211
rect 3801 3205 3803 3239
rect 3710 3203 3803 3205
rect 3817 3193 3821 3294
rect 4781 3295 4839 3298
rect 4351 3280 4376 3283
rect 4129 3274 4231 3277
rect 4129 3264 4132 3274
rect 4160 3264 4218 3267
rect 4094 3253 4137 3255
rect 4094 3197 4096 3253
rect 4109 3243 4111 3248
rect 4135 3243 4137 3253
rect 4160 3243 4162 3264
rect 4186 3243 4188 3247
rect 4109 3229 4111 3238
rect 4135 3235 4137 3238
rect 4109 3227 4137 3229
rect 4109 3212 4111 3215
rect 4135 3212 4137 3227
rect 4160 3226 4162 3238
rect 4160 3212 4162 3222
rect 4186 3212 4188 3238
rect 4196 3224 4202 3226
rect 4109 3197 4111 3207
rect 4094 3195 4111 3197
rect 3536 3176 3642 3179
rect 3717 3190 3821 3193
rect 4109 3190 4111 3195
rect 4135 3196 4137 3207
rect 4160 3204 4162 3207
rect 4135 3194 4141 3196
rect 4186 3196 4188 3207
rect 4145 3194 4188 3196
rect 4200 3190 4202 3224
rect 3312 3172 3314 3175
rect 3322 3172 3324 3175
rect 3182 3165 3184 3168
rect 3191 3165 3193 3168
rect 3182 3149 3184 3160
rect 3224 3165 3226 3168
rect 3154 3146 3184 3149
rect 3039 3139 3040 3143
rect 3006 3131 3007 3135
rect 3005 3128 3007 3131
rect 3038 3128 3040 3139
rect 3182 3134 3184 3146
rect 3191 3141 3193 3160
rect 3224 3149 3226 3160
rect 3192 3137 3193 3141
rect 3191 3134 3193 3137
rect 3224 3134 3226 3145
rect 2996 3120 2998 3123
rect 3005 3120 3007 3123
rect 3182 3126 3184 3129
rect 3191 3126 3193 3129
rect 3224 3126 3226 3129
rect 3038 3120 3040 3123
rect 3292 3106 3296 3152
rect 3312 3147 3314 3167
rect 3322 3156 3324 3167
rect 3368 3172 3370 3175
rect 3536 3167 3539 3176
rect 3312 3133 3314 3143
rect 3322 3133 3324 3152
rect 3368 3148 3370 3167
rect 3369 3144 3370 3148
rect 3536 3150 3539 3162
rect 3559 3166 3561 3169
rect 3568 3166 3570 3169
rect 3559 3150 3561 3161
rect 3601 3166 3603 3169
rect 3536 3147 3561 3150
rect 3368 3133 3370 3144
rect 3559 3135 3561 3147
rect 3568 3142 3570 3161
rect 3601 3150 3603 3161
rect 3717 3156 3720 3190
rect 4109 3188 4202 3190
rect 3875 3179 3877 3182
rect 3885 3179 3887 3182
rect 3745 3172 3747 3175
rect 3754 3172 3756 3175
rect 3745 3156 3747 3167
rect 3787 3172 3789 3175
rect 3717 3153 3747 3156
rect 3602 3146 3603 3150
rect 3569 3138 3570 3142
rect 3568 3135 3570 3138
rect 3601 3135 3603 3146
rect 3745 3141 3747 3153
rect 3754 3148 3756 3167
rect 3787 3156 3789 3167
rect 3755 3144 3756 3148
rect 3754 3141 3756 3144
rect 3787 3141 3789 3152
rect 3312 3125 3314 3128
rect 3322 3125 3324 3128
rect 3368 3125 3370 3128
rect 3559 3127 3561 3130
rect 3568 3127 3570 3130
rect 3745 3133 3747 3136
rect 3754 3133 3756 3136
rect 3787 3133 3789 3136
rect 3601 3127 3603 3130
rect 3855 3113 3859 3159
rect 3875 3154 3877 3174
rect 3885 3163 3887 3174
rect 3931 3179 3933 3182
rect 3875 3140 3877 3150
rect 3885 3140 3887 3159
rect 3931 3155 3933 3174
rect 4215 3165 4218 3264
rect 4302 3264 4305 3274
rect 4271 3254 4314 3256
rect 4271 3198 4273 3254
rect 4286 3244 4288 3249
rect 4312 3244 4314 3254
rect 4337 3244 4339 3247
rect 4286 3230 4288 3239
rect 4312 3236 4314 3239
rect 4337 3230 4339 3239
rect 4351 3230 4354 3280
rect 4715 3284 4758 3286
rect 4384 3280 4397 3283
rect 4363 3244 4365 3248
rect 4286 3228 4314 3230
rect 4286 3213 4288 3216
rect 4312 3213 4314 3228
rect 4337 3228 4354 3230
rect 4337 3227 4339 3228
rect 4337 3213 4339 3223
rect 4363 3213 4365 3239
rect 4373 3225 4379 3227
rect 4286 3198 4288 3208
rect 4271 3196 4288 3198
rect 4286 3191 4288 3196
rect 4312 3197 4314 3208
rect 4337 3205 4339 3208
rect 4312 3195 4334 3197
rect 4363 3197 4365 3208
rect 4338 3195 4365 3197
rect 4377 3191 4379 3225
rect 4286 3189 4379 3191
rect 4393 3179 4397 3280
rect 4715 3228 4717 3284
rect 4730 3274 4732 3279
rect 4756 3274 4758 3284
rect 4781 3274 4783 3295
rect 4807 3274 4809 3278
rect 4730 3260 4732 3269
rect 4756 3266 4758 3269
rect 4730 3258 4758 3260
rect 4730 3243 4732 3246
rect 4756 3243 4758 3258
rect 4781 3257 4783 3269
rect 4781 3243 4783 3253
rect 4807 3243 4809 3269
rect 4817 3255 4823 3257
rect 4730 3228 4732 3238
rect 4715 3226 4732 3228
rect 4730 3221 4732 3226
rect 4756 3227 4758 3238
rect 4781 3235 4783 3238
rect 4756 3225 4762 3227
rect 4807 3227 4809 3238
rect 4766 3225 4809 3227
rect 4821 3221 4823 3255
rect 4730 3219 4823 3221
rect 4836 3196 4839 3295
rect 4923 3295 4926 3313
rect 4972 3311 5020 3314
rect 4892 3285 4935 3287
rect 4892 3229 4894 3285
rect 4907 3275 4909 3280
rect 4933 3275 4935 3285
rect 4958 3275 4960 3278
rect 4907 3261 4909 3270
rect 4933 3267 4935 3270
rect 4958 3261 4960 3270
rect 4972 3261 4975 3311
rect 4984 3275 4986 3279
rect 4907 3259 4935 3261
rect 4907 3244 4909 3247
rect 4933 3244 4935 3259
rect 4958 3259 4975 3261
rect 4958 3258 4960 3259
rect 4958 3244 4960 3254
rect 4984 3244 4986 3270
rect 4994 3256 5000 3258
rect 4907 3229 4909 3239
rect 4892 3227 4909 3229
rect 4907 3222 4909 3227
rect 4933 3228 4935 3239
rect 4958 3236 4960 3239
rect 4933 3226 4955 3228
rect 4984 3228 4986 3239
rect 4959 3226 4986 3228
rect 4998 3222 5000 3256
rect 4907 3220 5000 3222
rect 5014 3210 5018 3311
rect 4725 3193 4839 3196
rect 4914 3207 5018 3210
rect 3932 3151 3933 3155
rect 3931 3140 3933 3151
rect 4110 3162 4218 3165
rect 4293 3176 4397 3179
rect 4110 3152 4113 3162
rect 4135 3152 4137 3155
rect 4144 3152 4146 3155
rect 3875 3132 3877 3135
rect 3885 3132 3887 3135
rect 4110 3136 4113 3146
rect 4135 3136 4137 3147
rect 4177 3152 4179 3155
rect 3931 3132 3933 3135
rect 4110 3133 4137 3136
rect 4135 3121 4137 3133
rect 4144 3128 4146 3147
rect 4177 3136 4179 3147
rect 4293 3142 4296 3176
rect 4451 3165 4453 3168
rect 4461 3165 4463 3168
rect 4321 3158 4323 3161
rect 4330 3158 4332 3161
rect 4321 3142 4323 3153
rect 4363 3158 4365 3161
rect 4293 3139 4323 3142
rect 4178 3132 4179 3136
rect 4145 3124 4146 3128
rect 4144 3121 4146 3124
rect 4177 3121 4179 3132
rect 4321 3127 4323 3139
rect 4330 3134 4332 3153
rect 4363 3142 4365 3153
rect 4331 3130 4332 3134
rect 4330 3127 4332 3130
rect 4363 3127 4365 3138
rect 4135 3113 4137 3116
rect 4144 3113 4146 3116
rect 4321 3119 4323 3122
rect 4330 3119 4332 3122
rect 4363 3119 4365 3122
rect 4177 3113 4179 3116
rect 3641 3109 3859 3113
rect 3078 3102 3296 3106
rect 4431 3099 4435 3145
rect 4451 3140 4453 3160
rect 4461 3149 4463 3160
rect 4507 3165 4509 3168
rect 4725 3167 4728 3186
rect 4756 3183 4758 3186
rect 4765 3183 4767 3186
rect 4756 3167 4758 3178
rect 4798 3183 4800 3186
rect 4725 3164 4758 3167
rect 4451 3126 4453 3136
rect 4461 3126 4463 3145
rect 4507 3141 4509 3160
rect 4756 3152 4758 3164
rect 4765 3159 4767 3178
rect 4798 3167 4800 3178
rect 4914 3173 4917 3207
rect 5072 3196 5074 3199
rect 5082 3196 5084 3199
rect 4942 3189 4944 3192
rect 4951 3189 4953 3192
rect 4942 3173 4944 3184
rect 4984 3189 4986 3192
rect 4914 3170 4944 3173
rect 4799 3163 4800 3167
rect 4766 3155 4767 3159
rect 4765 3152 4767 3155
rect 4798 3152 4800 3163
rect 4942 3158 4944 3170
rect 4951 3165 4953 3184
rect 4984 3173 4986 3184
rect 4952 3161 4953 3165
rect 4951 3158 4953 3161
rect 4984 3158 4986 3169
rect 4756 3144 4758 3147
rect 4765 3144 4767 3147
rect 4942 3150 4944 3153
rect 4951 3150 4953 3153
rect 4984 3150 4986 3153
rect 4798 3144 4800 3147
rect 4508 3137 4509 3141
rect 4507 3126 4509 3137
rect 4451 3118 4453 3121
rect 4461 3118 4463 3121
rect 5052 3130 5056 3176
rect 5072 3171 5074 3191
rect 5082 3180 5084 3191
rect 5128 3196 5130 3199
rect 5072 3157 5074 3167
rect 5082 3157 5084 3176
rect 5128 3172 5130 3191
rect 5129 3168 5130 3172
rect 5128 3157 5130 3168
rect 5072 3149 5074 3152
rect 5082 3149 5084 3152
rect 5128 3149 5130 3152
rect 4838 3126 5056 3130
rect 4507 3118 4509 3121
rect 4217 3095 4435 3099
rect 2950 3045 3172 3052
rect 1552 3008 2092 3013
rect 2335 3019 2789 3029
rect 242 2991 244 2994
rect 251 2991 253 2994
rect 242 2976 244 2986
rect 284 2991 286 2994
rect 243 2972 244 2976
rect 242 2960 244 2972
rect 251 2967 253 2986
rect 284 2975 286 2986
rect 285 2971 286 2975
rect 252 2963 253 2967
rect 251 2960 253 2963
rect 284 2960 286 2971
rect 242 2952 244 2955
rect 251 2952 253 2955
rect 284 2952 286 2955
rect 194 2949 228 2951
rect 179 2942 180 2945
rect 209 2941 231 2944
rect 194 2938 196 2941
rect 194 2924 196 2934
rect 227 2928 231 2941
rect 305 2932 309 2994
rect 1469 2981 1474 2983
rect 1469 2977 1755 2981
rect 1469 2932 1474 2977
rect 1866 2981 1950 2982
rect 1760 2978 1950 2981
rect 1760 2977 1865 2978
rect 2335 2982 2341 3019
rect 1955 2981 2089 2982
rect 2297 2981 2364 2982
rect 1955 2978 2163 2981
rect 2079 2977 2163 2978
rect 2168 2978 2364 2981
rect 2168 2977 2299 2978
rect 1774 2964 1776 2965
rect 1682 2950 1725 2952
rect 305 2929 1491 2932
rect 227 2925 269 2928
rect 190 2922 196 2924
rect 131 2918 173 2920
rect 131 2914 134 2918
rect 105 2907 107 2910
rect 114 2907 116 2910
rect 105 2892 107 2902
rect 147 2907 149 2910
rect 106 2888 107 2892
rect 105 2876 107 2888
rect 114 2883 116 2902
rect 147 2891 149 2902
rect 148 2887 149 2891
rect 115 2879 116 2883
rect 114 2876 116 2879
rect 147 2876 149 2887
rect 105 2868 107 2871
rect 114 2868 116 2871
rect 147 2868 149 2871
rect 58 2861 93 2864
rect 158 2825 161 2860
rect 170 2862 173 2918
rect 194 2915 196 2922
rect 266 2918 269 2925
rect 305 2917 309 2929
rect 426 2925 429 2929
rect 569 2925 572 2929
rect 731 2928 735 2929
rect 886 2928 891 2929
rect 732 2925 735 2928
rect 888 2925 891 2928
rect 1026 2925 1029 2929
rect 1169 2925 1172 2929
rect 1331 2928 1335 2929
rect 1469 2928 1474 2929
rect 1332 2925 1335 2928
rect 1488 2925 1491 2929
rect 301 2913 309 2917
rect 194 2908 196 2911
rect 241 2910 243 2913
rect 250 2910 252 2913
rect 206 2877 209 2903
rect 241 2895 243 2905
rect 283 2910 285 2913
rect 242 2891 243 2895
rect 241 2879 243 2891
rect 250 2886 252 2905
rect 283 2894 285 2905
rect 284 2890 285 2894
rect 251 2882 252 2886
rect 250 2879 252 2882
rect 283 2879 285 2890
rect 206 2874 233 2877
rect 230 2870 233 2874
rect 241 2871 243 2874
rect 250 2871 252 2874
rect 283 2871 285 2874
rect 170 2859 180 2862
rect 210 2859 235 2862
rect 194 2855 196 2858
rect 174 2825 177 2845
rect 194 2841 196 2851
rect 190 2839 196 2841
rect 194 2833 196 2839
rect 231 2836 235 2859
rect 305 2846 309 2913
rect 400 2917 402 2920
rect 409 2917 411 2920
rect 400 2902 402 2912
rect 442 2917 444 2920
rect 543 2917 545 2920
rect 552 2917 554 2920
rect 401 2898 402 2902
rect 400 2886 402 2898
rect 409 2893 411 2912
rect 442 2901 444 2912
rect 543 2902 545 2912
rect 585 2917 587 2920
rect 706 2917 708 2920
rect 715 2917 717 2920
rect 443 2897 444 2901
rect 544 2898 545 2902
rect 410 2889 411 2893
rect 409 2886 411 2889
rect 442 2886 444 2897
rect 400 2878 402 2881
rect 409 2878 411 2881
rect 543 2886 545 2898
rect 552 2893 554 2912
rect 585 2901 587 2912
rect 706 2902 708 2912
rect 748 2917 750 2920
rect 862 2917 864 2920
rect 871 2917 873 2920
rect 586 2897 587 2901
rect 707 2898 708 2902
rect 553 2889 554 2893
rect 552 2886 554 2889
rect 585 2886 587 2897
rect 442 2878 444 2881
rect 543 2878 545 2881
rect 552 2878 554 2881
rect 706 2886 708 2898
rect 715 2893 717 2912
rect 748 2901 750 2912
rect 862 2902 864 2912
rect 904 2917 906 2920
rect 1000 2917 1002 2920
rect 1009 2917 1011 2920
rect 749 2897 750 2901
rect 863 2898 864 2902
rect 716 2889 717 2893
rect 715 2886 717 2889
rect 748 2886 750 2897
rect 585 2878 587 2881
rect 706 2878 708 2881
rect 715 2878 717 2881
rect 862 2886 864 2898
rect 871 2893 873 2912
rect 904 2901 906 2912
rect 1000 2902 1002 2912
rect 1042 2917 1044 2920
rect 1143 2917 1145 2920
rect 1152 2917 1154 2920
rect 905 2897 906 2901
rect 1001 2898 1002 2902
rect 872 2889 873 2893
rect 871 2886 873 2889
rect 904 2886 906 2897
rect 748 2878 750 2881
rect 862 2878 864 2881
rect 871 2878 873 2881
rect 1000 2886 1002 2898
rect 1009 2893 1011 2912
rect 1042 2901 1044 2912
rect 1143 2902 1145 2912
rect 1185 2917 1187 2920
rect 1306 2917 1308 2920
rect 1315 2917 1317 2920
rect 1043 2897 1044 2901
rect 1144 2898 1145 2902
rect 1010 2889 1011 2893
rect 1009 2886 1011 2889
rect 1042 2886 1044 2897
rect 904 2878 906 2881
rect 1000 2878 1002 2881
rect 1009 2878 1011 2881
rect 1143 2886 1145 2898
rect 1152 2893 1154 2912
rect 1185 2901 1187 2912
rect 1306 2902 1308 2912
rect 1348 2917 1350 2920
rect 1462 2917 1464 2920
rect 1471 2917 1473 2920
rect 1186 2897 1187 2901
rect 1307 2898 1308 2902
rect 1153 2889 1154 2893
rect 1152 2886 1154 2889
rect 1185 2886 1187 2897
rect 1042 2878 1044 2881
rect 1143 2878 1145 2881
rect 1152 2878 1154 2881
rect 1306 2886 1308 2898
rect 1315 2893 1317 2912
rect 1348 2901 1350 2912
rect 1462 2902 1464 2912
rect 1504 2917 1506 2920
rect 1349 2897 1350 2901
rect 1463 2898 1464 2902
rect 1316 2889 1317 2893
rect 1315 2886 1317 2889
rect 1348 2886 1350 2897
rect 1185 2878 1187 2881
rect 1306 2878 1308 2881
rect 1315 2878 1317 2881
rect 1462 2886 1464 2898
rect 1471 2893 1473 2912
rect 1504 2901 1506 2912
rect 1505 2897 1506 2901
rect 1472 2889 1473 2893
rect 1471 2886 1473 2889
rect 1504 2886 1506 2897
rect 1348 2878 1350 2881
rect 1462 2878 1464 2881
rect 1471 2878 1473 2881
rect 1504 2878 1506 2881
rect 1626 2847 1631 2920
rect 1682 2894 1684 2950
rect 1697 2940 1699 2945
rect 1723 2940 1725 2950
rect 1748 2940 1750 2943
rect 1774 2940 1776 2958
rect 1877 2951 1920 2953
rect 1697 2926 1699 2935
rect 1723 2932 1725 2935
rect 1697 2924 1725 2926
rect 1697 2909 1699 2912
rect 1723 2909 1725 2924
rect 1748 2923 1750 2935
rect 1748 2909 1750 2919
rect 1774 2909 1776 2935
rect 1784 2921 1790 2923
rect 1697 2894 1699 2904
rect 1682 2892 1699 2894
rect 1697 2888 1699 2892
rect 1723 2893 1725 2904
rect 1748 2901 1750 2904
rect 1774 2893 1776 2904
rect 1723 2891 1776 2893
rect 1788 2888 1790 2921
rect 1877 2895 1879 2951
rect 1892 2941 1894 2946
rect 1918 2941 1920 2951
rect 1943 2941 1945 2946
rect 1969 2941 1971 2959
rect 2090 2950 2133 2952
rect 1892 2927 1894 2936
rect 1918 2933 1920 2936
rect 1892 2925 1920 2927
rect 1892 2910 1894 2913
rect 1918 2910 1920 2925
rect 1943 2924 1945 2936
rect 1943 2910 1945 2920
rect 1969 2910 1971 2936
rect 1979 2922 1985 2924
rect 1892 2895 1894 2905
rect 1877 2893 1894 2895
rect 1697 2886 1790 2888
rect 1892 2889 1894 2893
rect 1918 2894 1920 2905
rect 1943 2902 1945 2905
rect 1969 2894 1971 2905
rect 1918 2892 1971 2894
rect 1983 2889 1985 2922
rect 1892 2887 1985 2889
rect 2072 2857 2075 2900
rect 2090 2894 2092 2950
rect 2105 2940 2107 2945
rect 2131 2940 2133 2950
rect 2156 2940 2158 2944
rect 2182 2940 2184 2962
rect 2105 2926 2107 2935
rect 2131 2932 2133 2935
rect 2105 2924 2133 2926
rect 2105 2909 2107 2912
rect 2131 2909 2133 2924
rect 2156 2923 2158 2935
rect 2156 2909 2158 2919
rect 2182 2909 2184 2935
rect 2192 2921 2198 2923
rect 2105 2894 2107 2904
rect 2090 2892 2107 2894
rect 2105 2888 2107 2892
rect 2131 2893 2133 2904
rect 2156 2901 2158 2904
rect 2182 2893 2184 2904
rect 2131 2891 2184 2893
rect 2196 2888 2198 2921
rect 2105 2886 2198 2888
rect 2279 2847 2284 2964
rect 2291 2951 2334 2953
rect 2291 2895 2293 2951
rect 2306 2941 2308 2946
rect 2332 2941 2334 2951
rect 2357 2941 2359 2944
rect 2383 2941 2385 2986
rect 2306 2927 2308 2936
rect 2332 2933 2334 2936
rect 2306 2925 2334 2927
rect 2306 2910 2308 2913
rect 2332 2910 2334 2925
rect 2357 2924 2359 2936
rect 2357 2910 2359 2920
rect 2383 2910 2385 2936
rect 2393 2922 2399 2924
rect 2306 2895 2308 2905
rect 2291 2893 2308 2895
rect 2306 2889 2308 2893
rect 2332 2894 2334 2905
rect 2357 2902 2359 2905
rect 2383 2894 2385 2905
rect 2332 2892 2385 2894
rect 2397 2889 2399 2922
rect 2306 2887 2399 2889
rect 2950 2884 2957 3045
rect 3180 3045 3659 3052
rect 4843 3052 4850 3067
rect 3667 3045 4313 3052
rect 4321 3046 4850 3052
rect 4321 3045 4842 3046
rect 2648 2880 2958 2884
rect 305 2843 331 2846
rect 305 2840 309 2843
rect 231 2832 273 2836
rect 269 2831 273 2832
rect 194 2826 196 2829
rect 270 2827 273 2831
rect 158 2822 181 2825
rect 173 2598 177 2822
rect 306 2826 309 2840
rect 305 2822 309 2826
rect 205 2781 208 2821
rect 245 2819 247 2822
rect 254 2819 256 2822
rect 245 2804 247 2814
rect 287 2819 289 2822
rect 246 2800 247 2804
rect 245 2788 247 2800
rect 254 2795 256 2814
rect 287 2803 289 2814
rect 288 2799 289 2803
rect 255 2791 256 2795
rect 254 2788 256 2791
rect 287 2788 289 2799
rect 224 2783 237 2786
rect 224 2781 227 2783
rect 205 2778 227 2781
rect 234 2779 237 2783
rect 245 2780 247 2783
rect 254 2780 256 2783
rect 328 2783 331 2843
rect 1626 2841 2284 2847
rect 2109 2783 2171 2784
rect 287 2780 289 2783
rect 328 2780 2171 2783
rect 330 2658 334 2780
rect 426 2776 429 2780
rect 569 2776 572 2780
rect 731 2779 735 2780
rect 886 2779 891 2780
rect 732 2776 735 2779
rect 888 2776 891 2779
rect 1026 2776 1029 2780
rect 1169 2776 1172 2780
rect 1331 2779 1335 2780
rect 1332 2776 1335 2779
rect 1488 2776 1491 2780
rect 1607 2779 2171 2780
rect 400 2768 402 2771
rect 409 2768 411 2771
rect 400 2753 402 2763
rect 442 2768 444 2771
rect 543 2768 545 2771
rect 552 2768 554 2771
rect 401 2749 402 2753
rect 400 2737 402 2749
rect 409 2744 411 2763
rect 442 2752 444 2763
rect 543 2753 545 2763
rect 585 2768 587 2771
rect 706 2768 708 2771
rect 715 2768 717 2771
rect 443 2748 444 2752
rect 544 2749 545 2753
rect 410 2740 411 2744
rect 409 2737 411 2740
rect 442 2737 444 2748
rect 400 2729 402 2732
rect 409 2729 411 2732
rect 543 2737 545 2749
rect 552 2744 554 2763
rect 585 2752 587 2763
rect 706 2753 708 2763
rect 748 2768 750 2771
rect 862 2768 864 2771
rect 871 2768 873 2771
rect 586 2748 587 2752
rect 707 2749 708 2753
rect 553 2740 554 2744
rect 552 2737 554 2740
rect 585 2737 587 2748
rect 442 2729 444 2732
rect 543 2729 545 2732
rect 552 2729 554 2732
rect 706 2737 708 2749
rect 715 2744 717 2763
rect 748 2752 750 2763
rect 862 2753 864 2763
rect 904 2768 906 2771
rect 1000 2768 1002 2771
rect 1009 2768 1011 2771
rect 749 2748 750 2752
rect 863 2749 864 2753
rect 716 2740 717 2744
rect 715 2737 717 2740
rect 748 2737 750 2748
rect 585 2729 587 2732
rect 706 2729 708 2732
rect 715 2729 717 2732
rect 862 2737 864 2749
rect 871 2744 873 2763
rect 904 2752 906 2763
rect 1000 2753 1002 2763
rect 1042 2768 1044 2771
rect 1143 2768 1145 2771
rect 1152 2768 1154 2771
rect 905 2748 906 2752
rect 1001 2749 1002 2753
rect 872 2740 873 2744
rect 871 2737 873 2740
rect 904 2737 906 2748
rect 748 2729 750 2732
rect 862 2729 864 2732
rect 871 2729 873 2732
rect 1000 2737 1002 2749
rect 1009 2744 1011 2763
rect 1042 2752 1044 2763
rect 1143 2753 1145 2763
rect 1185 2768 1187 2771
rect 1306 2768 1308 2771
rect 1315 2768 1317 2771
rect 1043 2748 1044 2752
rect 1144 2749 1145 2753
rect 1010 2740 1011 2744
rect 1009 2737 1011 2740
rect 1042 2737 1044 2748
rect 904 2729 906 2732
rect 1000 2729 1002 2732
rect 1009 2729 1011 2732
rect 1143 2737 1145 2749
rect 1152 2744 1154 2763
rect 1185 2752 1187 2763
rect 1306 2753 1308 2763
rect 1348 2768 1350 2771
rect 1462 2768 1464 2771
rect 1471 2768 1473 2771
rect 1186 2748 1187 2752
rect 1307 2749 1308 2753
rect 1153 2740 1154 2744
rect 1152 2737 1154 2740
rect 1185 2737 1187 2748
rect 1042 2729 1044 2732
rect 1143 2729 1145 2732
rect 1152 2729 1154 2732
rect 1306 2737 1308 2749
rect 1315 2744 1317 2763
rect 1348 2752 1350 2763
rect 1462 2753 1464 2763
rect 1504 2768 1506 2771
rect 1349 2748 1350 2752
rect 1463 2749 1464 2753
rect 1316 2740 1317 2744
rect 1315 2737 1317 2740
rect 1348 2737 1350 2748
rect 1185 2729 1187 2732
rect 1306 2729 1308 2732
rect 1315 2729 1317 2732
rect 1462 2737 1464 2749
rect 1471 2744 1473 2763
rect 1504 2752 1506 2763
rect 1505 2748 1506 2752
rect 1472 2740 1473 2744
rect 1471 2737 1473 2740
rect 1504 2737 1506 2748
rect 1348 2729 1350 2732
rect 1462 2729 1464 2732
rect 1471 2729 1473 2732
rect 1504 2729 1506 2732
rect 2164 2703 2169 2779
rect 2369 2752 2371 2755
rect 2384 2752 2386 2755
rect 2399 2752 2401 2755
rect 2414 2752 2416 2755
rect 2428 2752 2430 2755
rect 2454 2752 2456 2755
rect 2369 2717 2371 2742
rect 2384 2717 2386 2742
rect 2399 2717 2401 2742
rect 2414 2717 2416 2742
rect 2428 2717 2430 2742
rect 2454 2726 2456 2742
rect 2471 2722 2711 2726
rect 2454 2717 2456 2722
rect 2123 2692 2125 2695
rect 2123 2675 2125 2688
rect 2369 2676 2371 2707
rect 2384 2688 2386 2707
rect 2399 2688 2401 2707
rect 2414 2688 2416 2707
rect 2428 2688 2430 2707
rect 2454 2704 2456 2707
rect 1987 2673 2125 2675
rect 330 2655 1491 2658
rect 426 2651 429 2655
rect 569 2651 572 2655
rect 400 2643 402 2646
rect 409 2643 411 2646
rect 400 2628 402 2638
rect 442 2643 444 2646
rect 543 2643 545 2646
rect 552 2643 554 2646
rect 401 2624 402 2628
rect 400 2612 402 2624
rect 409 2619 411 2638
rect 442 2627 444 2638
rect 543 2628 545 2638
rect 585 2643 587 2646
rect 443 2623 444 2627
rect 544 2624 545 2628
rect 410 2615 411 2619
rect 409 2612 411 2615
rect 442 2612 444 2623
rect 400 2604 402 2607
rect 409 2604 411 2607
rect 543 2612 545 2624
rect 552 2619 554 2638
rect 585 2627 587 2638
rect 586 2623 587 2627
rect 553 2615 554 2619
rect 552 2612 554 2615
rect 585 2612 587 2623
rect 442 2604 444 2607
rect 543 2604 545 2607
rect 552 2604 554 2607
rect 585 2604 587 2607
rect 173 2593 229 2598
rect 635 2299 639 2655
rect 731 2654 735 2655
rect 886 2654 891 2655
rect 732 2651 735 2654
rect 888 2651 891 2654
rect 1026 2651 1029 2655
rect 1169 2651 1172 2655
rect 1331 2654 1335 2655
rect 1332 2651 1335 2654
rect 1488 2651 1491 2655
rect 706 2643 708 2646
rect 715 2643 717 2646
rect 706 2628 708 2638
rect 748 2643 750 2646
rect 862 2643 864 2646
rect 871 2643 873 2646
rect 707 2624 708 2628
rect 706 2612 708 2624
rect 715 2619 717 2638
rect 748 2627 750 2638
rect 862 2628 864 2638
rect 904 2643 906 2646
rect 1000 2643 1002 2646
rect 1009 2643 1011 2646
rect 749 2623 750 2627
rect 863 2624 864 2628
rect 716 2615 717 2619
rect 715 2612 717 2615
rect 748 2612 750 2623
rect 706 2604 708 2607
rect 715 2604 717 2607
rect 862 2612 864 2624
rect 871 2619 873 2638
rect 904 2627 906 2638
rect 1000 2628 1002 2638
rect 1042 2643 1044 2646
rect 1143 2643 1145 2646
rect 1152 2643 1154 2646
rect 905 2623 906 2627
rect 1001 2624 1002 2628
rect 872 2615 873 2619
rect 871 2612 873 2615
rect 904 2612 906 2623
rect 748 2604 750 2607
rect 862 2604 864 2607
rect 871 2604 873 2607
rect 1000 2612 1002 2624
rect 1009 2619 1011 2638
rect 1042 2627 1044 2638
rect 1143 2628 1145 2638
rect 1185 2643 1187 2646
rect 1306 2643 1308 2646
rect 1315 2643 1317 2646
rect 1043 2623 1044 2627
rect 1144 2624 1145 2628
rect 1010 2615 1011 2619
rect 1009 2612 1011 2615
rect 1042 2612 1044 2623
rect 904 2604 906 2607
rect 1000 2604 1002 2607
rect 1009 2604 1011 2607
rect 1143 2612 1145 2624
rect 1152 2619 1154 2638
rect 1185 2627 1187 2638
rect 1306 2628 1308 2638
rect 1348 2643 1350 2646
rect 1462 2643 1464 2646
rect 1471 2643 1473 2646
rect 1186 2623 1187 2627
rect 1307 2624 1308 2628
rect 1153 2615 1154 2619
rect 1152 2612 1154 2615
rect 1185 2612 1187 2623
rect 1042 2604 1044 2607
rect 1143 2604 1145 2607
rect 1152 2604 1154 2607
rect 1306 2612 1308 2624
rect 1315 2619 1317 2638
rect 1348 2627 1350 2638
rect 1462 2628 1464 2638
rect 1504 2643 1506 2646
rect 1349 2623 1350 2627
rect 1463 2624 1464 2628
rect 1316 2615 1317 2619
rect 1315 2612 1317 2615
rect 1348 2612 1350 2623
rect 1185 2604 1187 2607
rect 1306 2604 1308 2607
rect 1315 2604 1317 2607
rect 1462 2612 1464 2624
rect 1471 2619 1473 2638
rect 1504 2627 1506 2638
rect 1505 2623 1506 2627
rect 1472 2615 1473 2619
rect 1471 2612 1473 2615
rect 1504 2612 1506 2623
rect 1348 2604 1350 2607
rect 1462 2604 1464 2607
rect 1471 2604 1473 2607
rect 1504 2604 1506 2607
rect 635 2296 1273 2299
rect 808 2292 811 2296
rect 951 2292 954 2296
rect 1113 2295 1117 2296
rect 1114 2292 1117 2295
rect 1270 2292 1273 2296
rect 782 2284 784 2287
rect 791 2284 793 2287
rect 782 2269 784 2279
rect 824 2284 826 2287
rect 925 2284 927 2287
rect 934 2284 936 2287
rect 783 2265 784 2269
rect 782 2253 784 2265
rect 791 2260 793 2279
rect 824 2268 826 2279
rect 925 2269 927 2279
rect 967 2284 969 2287
rect 1088 2284 1090 2287
rect 1097 2284 1099 2287
rect 825 2264 826 2268
rect 926 2265 927 2269
rect 792 2256 793 2260
rect 791 2253 793 2256
rect 824 2253 826 2264
rect 782 2245 784 2248
rect 791 2245 793 2248
rect 925 2253 927 2265
rect 934 2260 936 2279
rect 967 2268 969 2279
rect 1088 2269 1090 2279
rect 1130 2284 1132 2287
rect 1244 2284 1246 2287
rect 1253 2284 1255 2287
rect 968 2264 969 2268
rect 1089 2265 1090 2269
rect 935 2256 936 2260
rect 934 2253 936 2256
rect 967 2253 969 2264
rect 824 2245 826 2248
rect 925 2245 927 2248
rect 934 2245 936 2248
rect 1088 2253 1090 2265
rect 1097 2260 1099 2279
rect 1130 2268 1132 2279
rect 1244 2269 1246 2279
rect 1286 2284 1288 2287
rect 1131 2264 1132 2268
rect 1245 2265 1246 2269
rect 1098 2256 1099 2260
rect 1097 2253 1099 2256
rect 1130 2253 1132 2264
rect 967 2245 969 2248
rect 1088 2245 1090 2248
rect 1097 2245 1099 2248
rect 1244 2253 1246 2265
rect 1253 2260 1255 2279
rect 1286 2268 1288 2279
rect 1287 2264 1288 2268
rect 1254 2256 1255 2260
rect 1253 2253 1255 2256
rect 1286 2253 1288 2264
rect 1130 2245 1132 2248
rect 1244 2245 1246 2248
rect 1253 2245 1255 2248
rect 1286 2245 1288 2248
rect 1987 1841 1989 2673
rect 2123 2668 2125 2673
rect 2135 2672 2371 2676
rect 2123 2661 2125 2664
rect 2500 2652 2502 2655
rect 2515 2652 2517 2655
rect 2535 2652 2537 2655
rect 2545 2652 2547 2655
rect 2571 2652 2573 2655
rect 2708 2644 2711 2722
rect 2818 2699 2820 2702
rect 2830 2699 2832 2702
rect 2845 2699 2847 2702
rect 2855 2699 2857 2702
rect 2878 2699 2880 2702
rect 2818 2669 2820 2692
rect 2830 2669 2832 2692
rect 2845 2669 2847 2692
rect 2855 2669 2857 2692
rect 2878 2677 2880 2692
rect 2878 2669 2880 2673
rect 2818 2644 2820 2662
rect 2125 2626 2127 2629
rect 2125 2609 2127 2622
rect 2500 2617 2502 2642
rect 2515 2617 2517 2642
rect 2535 2617 2537 2642
rect 2545 2617 2547 2642
rect 2571 2626 2573 2642
rect 2708 2641 2820 2644
rect 2830 2626 2832 2662
rect 2588 2622 2832 2626
rect 2571 2617 2573 2622
rect 1994 2607 2127 2609
rect 1994 1989 1996 2607
rect 2125 2602 2127 2607
rect 2145 2606 2470 2610
rect 2638 2614 2640 2617
rect 2653 2614 2655 2617
rect 2673 2614 2675 2617
rect 2697 2614 2699 2617
rect 2125 2595 2127 2598
rect 2468 2588 2470 2606
rect 2500 2588 2502 2607
rect 2468 2586 2502 2588
rect 2128 2559 2130 2562
rect 2128 2542 2130 2555
rect 2001 2540 2130 2542
rect 2001 2143 2003 2540
rect 2128 2535 2130 2540
rect 2128 2528 2130 2531
rect 2128 2492 2130 2495
rect 2128 2475 2130 2488
rect 2018 2473 2130 2475
rect 2018 2304 2020 2473
rect 2128 2468 2130 2473
rect 2128 2461 2130 2464
rect 2146 2387 2148 2390
rect 2031 2380 2067 2382
rect 2018 2301 2023 2304
rect 2031 2295 2033 2380
rect 2046 2351 2048 2354
rect 2065 2351 2067 2380
rect 2146 2370 2148 2383
rect 2141 2368 2148 2370
rect 2146 2363 2148 2368
rect 2146 2356 2148 2359
rect 2090 2351 2092 2354
rect 2109 2351 2111 2354
rect 2046 2334 2048 2346
rect 2065 2343 2067 2346
rect 2090 2334 2092 2346
rect 2046 2332 2067 2334
rect 2046 2320 2048 2323
rect 2065 2320 2067 2332
rect 2091 2330 2092 2334
rect 2090 2320 2092 2330
rect 2109 2320 2111 2346
rect 2120 2331 2126 2333
rect 2046 2295 2048 2315
rect 2065 2304 2067 2315
rect 2090 2312 2092 2315
rect 2109 2304 2111 2315
rect 2069 2302 2111 2304
rect 2124 2295 2126 2331
rect 2031 2293 2126 2295
rect 2148 2226 2150 2229
rect 2033 2219 2069 2221
rect 2001 2140 2025 2143
rect 2033 2134 2035 2219
rect 2048 2190 2050 2193
rect 2067 2190 2069 2219
rect 2148 2209 2150 2222
rect 2143 2207 2150 2209
rect 2148 2202 2150 2207
rect 2148 2195 2150 2198
rect 2092 2190 2094 2193
rect 2111 2190 2113 2193
rect 2048 2173 2050 2185
rect 2067 2182 2069 2185
rect 2092 2173 2094 2185
rect 2048 2171 2069 2173
rect 2048 2159 2050 2162
rect 2067 2159 2069 2171
rect 2093 2169 2094 2173
rect 2092 2159 2094 2169
rect 2111 2159 2113 2185
rect 2122 2170 2128 2172
rect 2048 2134 2050 2154
rect 2067 2143 2069 2154
rect 2092 2151 2094 2154
rect 2111 2143 2113 2154
rect 2071 2141 2113 2143
rect 2126 2134 2128 2170
rect 2033 2132 2128 2134
rect 2515 2095 2517 2607
rect 2535 2588 2537 2607
rect 2545 2587 2547 2607
rect 2571 2604 2573 2607
rect 2638 2579 2640 2604
rect 2653 2579 2655 2604
rect 2673 2579 2675 2604
rect 2697 2588 2699 2604
rect 2845 2588 2847 2662
rect 2714 2584 2847 2588
rect 2697 2579 2699 2584
rect 2764 2569 2766 2572
rect 2785 2569 2787 2572
rect 2811 2569 2813 2572
rect 2638 2550 2640 2569
rect 2653 2528 2655 2569
rect 2673 2549 2675 2569
rect 2697 2566 2699 2569
rect 2764 2541 2766 2564
rect 2785 2541 2787 2564
rect 2811 2552 2813 2565
rect 2855 2553 2857 2662
rect 2878 2659 2880 2662
rect 2806 2550 2813 2552
rect 2811 2545 2813 2550
rect 2822 2549 2857 2553
rect 2811 2538 2813 2541
rect 2764 2476 2766 2534
rect 2785 2523 2787 2534
rect 2578 2472 2766 2476
rect 2917 2284 2962 2289
rect 2747 2178 2749 2181
rect 2762 2178 2764 2181
rect 2782 2178 2784 2181
rect 2792 2178 2794 2181
rect 2818 2178 2820 2181
rect 2747 2143 2749 2168
rect 2762 2143 2764 2168
rect 2782 2143 2784 2168
rect 2792 2143 2794 2168
rect 2818 2152 2820 2168
rect 2906 2169 2908 2172
rect 2917 2169 2919 2284
rect 2906 2152 2908 2164
rect 2948 2169 2950 2172
rect 2818 2143 2820 2148
rect 2906 2138 2908 2147
rect 2917 2138 2919 2164
rect 2948 2153 2950 2164
rect 2949 2149 2950 2153
rect 2948 2138 2950 2149
rect 2747 2116 2749 2133
rect 2724 2114 2749 2116
rect 2762 2109 2764 2133
rect 2724 2107 2764 2109
rect 2782 2101 2784 2133
rect 2724 2099 2784 2101
rect 2062 2091 2517 2095
rect 2792 2093 2794 2133
rect 2818 2130 2820 2133
rect 2906 2130 2908 2133
rect 2917 2130 2919 2133
rect 2948 2130 2950 2133
rect 2724 2091 2794 2093
rect 2147 2072 2149 2075
rect 2032 2065 2068 2067
rect 1994 1986 2024 1989
rect 2032 1980 2034 2065
rect 2047 2036 2049 2039
rect 2066 2036 2068 2065
rect 2147 2055 2149 2068
rect 2142 2053 2149 2055
rect 2147 2048 2149 2053
rect 2147 2041 2149 2044
rect 2091 2036 2093 2039
rect 2110 2036 2112 2039
rect 2047 2019 2049 2031
rect 2066 2028 2068 2031
rect 2091 2019 2093 2031
rect 2047 2017 2068 2019
rect 2047 2005 2049 2008
rect 2066 2005 2068 2017
rect 2092 2015 2093 2019
rect 2091 2005 2093 2015
rect 2110 2005 2112 2031
rect 2121 2016 2127 2018
rect 2047 1980 2049 2000
rect 2066 1989 2068 2000
rect 2091 1997 2093 2000
rect 2110 1989 2112 2000
rect 2070 1987 2112 1989
rect 2125 1980 2127 2016
rect 2032 1978 2127 1980
rect 2147 1924 2149 1927
rect 2032 1917 2068 1919
rect 1987 1838 2024 1841
rect 2032 1832 2034 1917
rect 2047 1888 2049 1891
rect 2066 1888 2068 1917
rect 2147 1907 2149 1920
rect 2809 1919 2811 1922
rect 2821 1919 2823 1922
rect 2836 1919 2838 1922
rect 2846 1919 2848 1922
rect 2869 1919 2871 1922
rect 2142 1905 2149 1907
rect 2147 1900 2149 1905
rect 2147 1893 2149 1896
rect 2091 1888 2093 1891
rect 2110 1888 2112 1891
rect 2809 1889 2811 1912
rect 2821 1889 2823 1912
rect 2836 1889 2838 1912
rect 2846 1889 2848 1912
rect 2869 1897 2871 1912
rect 2869 1889 2871 1893
rect 2047 1871 2049 1883
rect 2066 1880 2068 1883
rect 2091 1871 2093 1883
rect 2047 1869 2068 1871
rect 2047 1857 2049 1860
rect 2066 1857 2068 1869
rect 2092 1867 2093 1871
rect 2091 1857 2093 1867
rect 2110 1857 2112 1883
rect 2121 1868 2127 1870
rect 2047 1832 2049 1852
rect 2066 1841 2068 1852
rect 2091 1849 2093 1852
rect 2110 1841 2112 1852
rect 2070 1839 2112 1841
rect 2125 1832 2127 1868
rect 2584 1863 2586 1866
rect 2599 1863 2601 1866
rect 2614 1863 2616 1866
rect 2629 1863 2631 1866
rect 2643 1863 2645 1866
rect 2669 1863 2671 1866
rect 2032 1830 2127 1832
rect 2584 1828 2586 1853
rect 2599 1828 2601 1853
rect 2614 1828 2616 1853
rect 2629 1828 2631 1853
rect 2643 1828 2645 1853
rect 2669 1837 2671 1853
rect 2809 1837 2811 1882
rect 2686 1833 2811 1837
rect 2669 1828 2671 1833
rect 2123 1797 2125 1800
rect 2584 1798 2586 1818
rect 2599 1798 2601 1818
rect 2614 1798 2616 1818
rect 2629 1799 2631 1818
rect 2643 1799 2645 1818
rect 2669 1815 2671 1818
rect 2362 1795 2586 1798
rect 2123 1780 2125 1793
rect 2362 1781 2367 1795
rect 2105 1778 2125 1780
rect 2123 1773 2125 1778
rect 2189 1777 2367 1781
rect 2452 1779 2454 1782
rect 2467 1779 2469 1782
rect 2487 1779 2489 1782
rect 2497 1779 2499 1782
rect 2523 1779 2525 1782
rect 2123 1766 2125 1769
rect 2452 1744 2454 1769
rect 2467 1744 2469 1769
rect 2487 1744 2489 1769
rect 2497 1744 2499 1769
rect 2523 1753 2525 1769
rect 2821 1753 2823 1882
rect 2836 1869 2838 1882
rect 2540 1749 2823 1753
rect 2523 1744 2525 1749
rect 2125 1731 2127 1734
rect 2125 1714 2127 1727
rect 2452 1715 2454 1734
rect 2467 1715 2469 1734
rect 2487 1716 2489 1734
rect 2497 1716 2499 1734
rect 2523 1731 2525 1734
rect 2105 1712 2127 1714
rect 2125 1707 2127 1712
rect 2146 1712 2454 1715
rect 2311 1704 2313 1707
rect 2326 1704 2328 1707
rect 2346 1704 2348 1707
rect 2370 1704 2372 1707
rect 2125 1700 2127 1703
rect 2311 1669 2313 1694
rect 2326 1669 2328 1694
rect 2346 1669 2348 1694
rect 2370 1678 2372 1694
rect 2370 1669 2372 1674
rect 2128 1664 2130 1667
rect 2128 1647 2130 1660
rect 2105 1645 2130 1647
rect 2128 1640 2130 1645
rect 2140 1644 2293 1648
rect 2290 1638 2293 1644
rect 2311 1638 2313 1659
rect 2326 1640 2328 1659
rect 2128 1633 2130 1636
rect 2290 1635 2313 1638
rect 2346 1639 2348 1659
rect 2370 1656 2372 1659
rect 2213 1625 2215 1628
rect 2234 1625 2236 1628
rect 2260 1625 2262 1628
rect 2128 1597 2130 1600
rect 2213 1597 2215 1620
rect 2234 1597 2236 1620
rect 2260 1608 2262 1621
rect 2846 1609 2848 1882
rect 2869 1879 2871 1882
rect 2255 1606 2262 1608
rect 2260 1601 2262 1606
rect 2271 1605 2848 1609
rect 2128 1580 2130 1593
rect 2260 1594 2262 1597
rect 2213 1581 2215 1590
rect 2105 1578 2130 1580
rect 2128 1573 2130 1578
rect 2141 1577 2215 1581
rect 2234 1577 2236 1590
rect 2128 1566 2130 1569
<< polycontact >>
rect 208 3721 220 3733
rect 794 3639 804 3649
rect 1984 3648 1992 3657
rect 1335 3618 1343 3626
rect 2095 3605 2099 3609
rect 335 3581 339 3585
rect 232 3566 236 3571
rect 262 3529 266 3533
rect 296 3530 300 3534
rect 245 3501 249 3505
rect 406 3567 410 3571
rect 475 3586 482 3593
rect 439 3530 443 3534
rect 473 3531 477 3535
rect 438 3502 442 3506
rect 898 3588 902 3592
rect 795 3573 799 3578
rect 825 3536 829 3540
rect 859 3537 863 3541
rect 808 3508 812 3512
rect 217 3458 222 3464
rect 969 3574 973 3578
rect 1033 3593 1039 3598
rect 1002 3537 1006 3541
rect 1036 3538 1040 3542
rect 1001 3509 1005 3513
rect 1992 3590 1996 3595
rect 1474 3574 1478 3578
rect 1371 3559 1375 3564
rect 1401 3522 1405 3526
rect 1435 3523 1439 3527
rect 1384 3494 1388 3498
rect 278 3439 282 3443
rect 245 3431 249 3435
rect 464 3445 469 3449
rect 431 3437 435 3441
rect 535 3452 540 3456
rect 314 3401 321 3407
rect 562 3452 567 3456
rect 552 3443 557 3447
rect 778 3462 782 3467
rect 608 3444 612 3448
rect 841 3446 845 3450
rect 808 3438 812 3442
rect 1027 3452 1032 3456
rect 994 3444 998 3448
rect 1098 3459 1103 3463
rect 877 3408 884 3414
rect 1125 3459 1130 3463
rect 1115 3450 1120 3454
rect 1545 3560 1549 3564
rect 1619 3578 1627 3586
rect 1578 3523 1582 3527
rect 1612 3524 1616 3528
rect 1577 3495 1581 3499
rect 2022 3553 2026 3557
rect 2056 3554 2060 3558
rect 2005 3525 2009 3529
rect 2166 3591 2170 3595
rect 2199 3554 2203 3558
rect 2233 3555 2237 3559
rect 2256 3557 2264 3564
rect 2198 3526 2202 3530
rect 1964 3486 1972 3493
rect 1171 3451 1175 3455
rect 1353 3446 1359 3452
rect 1417 3432 1421 3436
rect 1384 3424 1388 3428
rect 1603 3438 1608 3442
rect 1570 3430 1574 3434
rect 1674 3445 1679 3449
rect 1453 3394 1460 3400
rect 1701 3445 1706 3449
rect 1691 3436 1696 3440
rect 2038 3463 2042 3467
rect 2005 3455 2009 3459
rect 2224 3469 2229 3473
rect 2191 3461 2195 3465
rect 2295 3476 2300 3480
rect 1747 3437 1751 3441
rect 2074 3425 2081 3431
rect 2322 3476 2327 3480
rect 2312 3467 2317 3471
rect 2368 3468 2372 3472
rect 2965 3421 2977 3433
rect 2085 3367 2095 3374
rect 415 3344 423 3353
rect 902 3345 910 3353
rect 1556 3344 1564 3352
rect 169 2948 173 2952
rect 426 3063 430 3067
rect 569 3063 573 3067
rect 732 3063 736 3067
rect 888 3063 892 3067
rect 1026 3063 1030 3067
rect 1169 3063 1173 3067
rect 1332 3063 1336 3067
rect 1488 3063 1492 3067
rect 397 3040 401 3044
rect 439 3039 443 3043
rect 540 3040 544 3044
rect 406 3031 410 3035
rect 582 3039 586 3043
rect 703 3040 707 3044
rect 549 3031 553 3035
rect 745 3039 749 3043
rect 859 3040 863 3044
rect 712 3031 716 3035
rect 901 3039 905 3043
rect 997 3040 1001 3044
rect 868 3031 872 3035
rect 1039 3039 1043 3043
rect 1140 3040 1144 3044
rect 1006 3031 1010 3035
rect 1182 3039 1186 3043
rect 1303 3040 1307 3044
rect 1149 3031 1153 3035
rect 1345 3039 1349 3043
rect 1459 3040 1463 3044
rect 1312 3031 1316 3035
rect 1501 3039 1505 3043
rect 1468 3031 1472 3035
rect 1541 3005 1552 3014
rect 3551 3339 3561 3349
rect 5013 3388 5023 3396
rect 4741 3348 4749 3357
rect 4092 3318 4100 3326
rect 4852 3305 4856 3309
rect 3092 3281 3096 3285
rect 2989 3266 2993 3271
rect 3019 3229 3023 3233
rect 3053 3230 3057 3234
rect 3002 3201 3006 3205
rect 3163 3267 3167 3271
rect 3232 3286 3239 3293
rect 3196 3230 3200 3234
rect 3230 3231 3234 3235
rect 3195 3202 3199 3206
rect 3655 3288 3659 3292
rect 3552 3273 3556 3278
rect 3582 3236 3586 3240
rect 3616 3237 3620 3241
rect 3565 3208 3569 3212
rect 2974 3158 2979 3164
rect 3726 3274 3730 3278
rect 3790 3293 3796 3298
rect 3759 3237 3763 3241
rect 3793 3238 3797 3242
rect 3758 3209 3762 3213
rect 4749 3290 4753 3295
rect 4231 3274 4235 3278
rect 4128 3259 4132 3264
rect 4158 3222 4162 3226
rect 4192 3223 4196 3227
rect 4141 3194 4145 3198
rect 3035 3139 3039 3143
rect 3002 3131 3006 3135
rect 3221 3145 3226 3149
rect 3188 3137 3192 3141
rect 3292 3152 3297 3156
rect 3071 3101 3078 3107
rect 3319 3152 3324 3156
rect 3309 3143 3314 3147
rect 3535 3162 3539 3167
rect 3365 3144 3369 3148
rect 3598 3146 3602 3150
rect 3565 3138 3569 3142
rect 3784 3152 3789 3156
rect 3751 3144 3755 3148
rect 3855 3159 3860 3163
rect 3634 3108 3641 3114
rect 3882 3159 3887 3163
rect 3872 3150 3877 3154
rect 4302 3260 4306 3264
rect 4376 3278 4384 3286
rect 4335 3223 4339 3227
rect 4369 3224 4373 3228
rect 4334 3195 4338 3199
rect 4779 3253 4783 3257
rect 4813 3254 4817 3258
rect 4762 3225 4766 3229
rect 4923 3291 4927 3295
rect 4956 3254 4960 3258
rect 4990 3255 4994 3259
rect 4955 3226 4959 3230
rect 4721 3186 4729 3193
rect 3928 3151 3932 3155
rect 4110 3146 4116 3152
rect 4174 3132 4178 3136
rect 4141 3124 4145 3128
rect 4360 3138 4365 3142
rect 4327 3130 4331 3134
rect 4431 3145 4436 3149
rect 4210 3094 4217 3100
rect 4458 3145 4463 3149
rect 4448 3136 4453 3140
rect 4795 3163 4799 3167
rect 4762 3155 4766 3159
rect 4981 3169 4986 3173
rect 4948 3161 4952 3165
rect 5052 3176 5057 3180
rect 4504 3137 4508 3141
rect 4831 3125 4838 3131
rect 5079 3176 5084 3180
rect 5069 3167 5074 3171
rect 5125 3168 5129 3172
rect 4842 3067 4852 3074
rect 268 2995 272 2999
rect 305 2994 309 3000
rect 239 2972 243 2976
rect 281 2971 285 2975
rect 248 2963 252 2967
rect 190 2948 194 2952
rect 228 2948 232 2952
rect 180 2941 184 2945
rect 205 2941 209 2945
rect 186 2921 190 2925
rect 1755 2976 1760 2982
rect 1950 2977 1955 2983
rect 2381 2986 2387 2992
rect 2163 2976 2168 2981
rect 2364 2977 2369 2983
rect 1772 2958 1779 2964
rect 1968 2959 1974 2965
rect 2181 2962 2186 2967
rect 2277 2964 2284 2970
rect 131 2910 135 2914
rect 102 2888 106 2892
rect 144 2887 148 2891
rect 111 2879 115 2883
rect 93 2860 97 2864
rect 157 2860 161 2864
rect 266 2914 270 2918
rect 426 2921 430 2925
rect 569 2921 573 2925
rect 732 2921 736 2925
rect 888 2921 892 2925
rect 1026 2921 1030 2925
rect 1169 2921 1173 2925
rect 1332 2921 1336 2925
rect 1488 2921 1492 2925
rect 1624 2920 1632 2927
rect 297 2913 301 2917
rect 205 2903 209 2907
rect 238 2891 242 2895
rect 280 2890 284 2894
rect 247 2882 251 2886
rect 230 2866 234 2870
rect 180 2858 184 2862
rect 206 2858 210 2862
rect 173 2845 177 2849
rect 186 2838 190 2842
rect 397 2898 401 2902
rect 439 2897 443 2901
rect 540 2898 544 2902
rect 406 2889 410 2893
rect 582 2897 586 2901
rect 703 2898 707 2902
rect 549 2889 553 2893
rect 745 2897 749 2901
rect 859 2898 863 2902
rect 712 2889 716 2893
rect 901 2897 905 2901
rect 997 2898 1001 2902
rect 868 2889 872 2893
rect 1039 2897 1043 2901
rect 1140 2898 1144 2902
rect 1006 2889 1010 2893
rect 1182 2897 1186 2901
rect 1303 2898 1307 2902
rect 1149 2889 1153 2893
rect 1345 2897 1349 2901
rect 1459 2898 1463 2902
rect 1312 2889 1316 2893
rect 1501 2897 1505 2901
rect 1468 2889 1472 2893
rect 1746 2919 1750 2923
rect 1780 2920 1784 2924
rect 1941 2920 1945 2924
rect 1975 2921 1979 2925
rect 2070 2900 2077 2907
rect 2154 2919 2158 2923
rect 2188 2920 2192 2924
rect 2071 2851 2077 2857
rect 2355 2920 2359 2924
rect 2389 2921 2393 2925
rect 2636 2877 2648 2887
rect 3172 3044 3180 3053
rect 3659 3045 3667 3053
rect 4313 3044 4321 3052
rect 181 2821 185 2825
rect 204 2821 208 2825
rect 270 2823 274 2827
rect 301 2822 305 2826
rect 242 2800 246 2804
rect 284 2799 288 2803
rect 251 2791 255 2795
rect 234 2775 238 2779
rect 426 2772 430 2776
rect 569 2772 573 2776
rect 732 2772 736 2776
rect 888 2772 892 2776
rect 1026 2772 1030 2776
rect 1169 2772 1173 2776
rect 1332 2772 1336 2776
rect 1488 2772 1492 2776
rect 397 2749 401 2753
rect 439 2748 443 2752
rect 540 2749 544 2753
rect 406 2740 410 2744
rect 582 2748 586 2752
rect 703 2749 707 2753
rect 549 2740 553 2744
rect 745 2748 749 2752
rect 859 2749 863 2753
rect 712 2740 716 2744
rect 901 2748 905 2752
rect 997 2749 1001 2753
rect 868 2740 872 2744
rect 1039 2748 1043 2752
rect 1140 2749 1144 2753
rect 1006 2740 1010 2744
rect 1182 2748 1186 2752
rect 1303 2749 1307 2753
rect 1149 2740 1153 2744
rect 1345 2748 1349 2752
rect 1459 2749 1463 2753
rect 1312 2740 1316 2744
rect 1501 2748 1505 2752
rect 1468 2740 1472 2744
rect 2452 2722 2456 2726
rect 2467 2722 2471 2726
rect 2164 2696 2172 2703
rect 2383 2684 2387 2688
rect 2398 2684 2402 2688
rect 2413 2684 2417 2688
rect 2427 2684 2431 2688
rect 426 2647 430 2651
rect 569 2647 573 2651
rect 397 2624 401 2628
rect 439 2623 443 2627
rect 540 2624 544 2628
rect 406 2615 410 2619
rect 582 2623 586 2627
rect 549 2615 553 2619
rect 229 2591 239 2599
rect 732 2647 736 2651
rect 888 2647 892 2651
rect 1026 2647 1030 2651
rect 1169 2647 1173 2651
rect 1332 2647 1336 2651
rect 1488 2647 1492 2651
rect 703 2624 707 2628
rect 745 2623 749 2627
rect 859 2624 863 2628
rect 712 2615 716 2619
rect 901 2623 905 2627
rect 997 2624 1001 2628
rect 868 2615 872 2619
rect 1039 2623 1043 2627
rect 1140 2624 1144 2628
rect 1006 2615 1010 2619
rect 1182 2623 1186 2627
rect 1303 2624 1307 2628
rect 1149 2615 1153 2619
rect 1345 2623 1349 2627
rect 1459 2624 1463 2628
rect 1312 2615 1316 2619
rect 1501 2623 1505 2627
rect 1468 2615 1472 2619
rect 808 2288 812 2292
rect 951 2288 955 2292
rect 1114 2288 1118 2292
rect 1270 2288 1274 2292
rect 779 2265 783 2269
rect 821 2264 825 2268
rect 922 2265 926 2269
rect 788 2256 792 2260
rect 964 2264 968 2268
rect 1085 2265 1089 2269
rect 931 2256 935 2260
rect 1127 2264 1131 2268
rect 1241 2265 1245 2269
rect 1094 2256 1098 2260
rect 1283 2264 1287 2268
rect 1250 2256 1254 2260
rect 2131 2672 2135 2676
rect 2876 2673 2880 2677
rect 2569 2622 2573 2626
rect 2584 2622 2588 2626
rect 2141 2606 2145 2610
rect 2023 2300 2027 2304
rect 2137 2367 2141 2371
rect 2087 2330 2091 2334
rect 2116 2330 2120 2334
rect 2065 2300 2069 2304
rect 2025 2139 2029 2143
rect 2139 2206 2143 2210
rect 2089 2169 2093 2173
rect 2118 2169 2122 2173
rect 2067 2139 2071 2143
rect 2534 2584 2538 2588
rect 2544 2583 2548 2587
rect 2695 2584 2699 2588
rect 2710 2584 2714 2588
rect 2637 2546 2641 2550
rect 2672 2545 2676 2549
rect 2802 2549 2806 2553
rect 2818 2549 2822 2553
rect 2652 2524 2656 2528
rect 2784 2519 2788 2523
rect 2574 2472 2578 2476
rect 2962 2282 2971 2292
rect 2816 2148 2820 2152
rect 2904 2147 2908 2152
rect 2945 2149 2949 2153
rect 2720 2114 2724 2118
rect 2720 2106 2724 2110
rect 2720 2098 2724 2102
rect 2058 2091 2062 2095
rect 2720 2090 2724 2094
rect 2024 1985 2028 1989
rect 2138 2052 2142 2056
rect 2088 2015 2092 2019
rect 2117 2015 2121 2019
rect 2066 1985 2070 1989
rect 2024 1837 2028 1841
rect 2138 1904 2142 1908
rect 2867 1893 2871 1897
rect 2088 1867 2092 1871
rect 2117 1867 2121 1871
rect 2066 1837 2070 1841
rect 2667 1833 2671 1837
rect 2682 1833 2686 1837
rect 2101 1777 2105 1781
rect 2598 1794 2602 1798
rect 2613 1794 2617 1798
rect 2628 1795 2632 1799
rect 2642 1795 2646 1799
rect 2185 1777 2189 1781
rect 2835 1865 2839 1869
rect 2521 1749 2525 1753
rect 2536 1749 2540 1753
rect 2101 1711 2105 1715
rect 2142 1711 2146 1715
rect 2466 1711 2470 1715
rect 2486 1712 2490 1716
rect 2496 1712 2500 1716
rect 2368 1674 2372 1678
rect 2101 1644 2105 1648
rect 2136 1644 2140 1648
rect 2325 1636 2329 1640
rect 2345 1635 2349 1639
rect 2251 1605 2255 1609
rect 2267 1605 2271 1609
rect 2101 1577 2105 1581
rect 2137 1577 2141 1581
rect 2233 1573 2237 1577
<< metal1 >>
rect 210 3616 215 3721
rect 1544 3670 2448 3676
rect 405 3663 411 3664
rect 400 3657 1222 3663
rect 405 3634 411 3657
rect 968 3639 973 3640
rect 404 3628 481 3634
rect 475 3593 481 3628
rect 794 3619 802 3639
rect 966 3634 1366 3639
rect 968 3628 973 3634
rect 968 3623 1038 3628
rect 1034 3598 1038 3623
rect 1544 3619 1550 3670
rect 1573 3634 1574 3639
rect 1583 3634 1789 3639
rect 1986 3638 1991 3648
rect 208 3574 255 3578
rect 208 3549 212 3574
rect 208 3519 212 3545
rect 217 3566 232 3570
rect 236 3566 247 3570
rect 217 3549 221 3566
rect 243 3549 247 3566
rect 217 3519 221 3545
rect 234 3519 238 3545
rect 243 3519 247 3545
rect 251 3533 255 3574
rect 259 3561 276 3565
rect 282 3561 288 3565
rect 259 3550 263 3561
rect 284 3551 288 3561
rect 251 3529 262 3533
rect 269 3525 273 3545
rect 251 3521 273 3525
rect 234 3512 238 3515
rect 251 3512 255 3521
rect 269 3519 273 3521
rect 234 3508 255 3512
rect 293 3534 297 3545
rect 293 3530 296 3534
rect 293 3519 297 3530
rect 259 3510 262 3514
rect 259 3507 277 3510
rect 285 3510 288 3514
rect 282 3507 288 3510
rect 245 3481 248 3501
rect 335 3491 339 3581
rect 771 3581 818 3585
rect 385 3575 432 3579
rect 385 3550 389 3575
rect 385 3520 389 3546
rect 394 3567 406 3571
rect 410 3567 424 3571
rect 394 3550 398 3567
rect 420 3550 424 3567
rect 394 3520 398 3546
rect 411 3520 415 3546
rect 420 3520 424 3546
rect 428 3534 432 3575
rect 436 3562 442 3566
rect 448 3562 465 3566
rect 436 3551 440 3562
rect 461 3552 465 3562
rect 771 3556 775 3581
rect 428 3530 439 3534
rect 446 3526 450 3546
rect 428 3522 450 3526
rect 411 3513 415 3516
rect 428 3513 432 3522
rect 446 3520 450 3522
rect 411 3509 432 3513
rect 470 3535 474 3546
rect 470 3531 473 3535
rect 470 3520 474 3531
rect 771 3526 775 3552
rect 780 3573 795 3577
rect 799 3573 810 3577
rect 780 3556 784 3573
rect 806 3556 810 3573
rect 780 3526 784 3552
rect 797 3526 801 3552
rect 806 3526 810 3552
rect 814 3540 818 3581
rect 822 3568 839 3572
rect 845 3568 851 3572
rect 822 3557 826 3568
rect 847 3558 851 3568
rect 814 3536 825 3540
rect 832 3532 836 3552
rect 814 3528 836 3532
rect 436 3512 440 3515
rect 797 3519 801 3522
rect 814 3519 818 3528
rect 832 3526 836 3528
rect 797 3515 818 3519
rect 856 3541 860 3552
rect 856 3537 859 3541
rect 856 3526 860 3537
rect 822 3517 825 3521
rect 436 3509 448 3512
rect 461 3512 465 3515
rect 822 3514 840 3517
rect 848 3517 851 3521
rect 845 3514 851 3517
rect 453 3509 465 3512
rect 438 3491 441 3502
rect 335 3488 441 3491
rect 808 3488 811 3508
rect 898 3498 902 3588
rect 948 3582 995 3586
rect 948 3557 952 3582
rect 948 3527 952 3553
rect 957 3574 969 3578
rect 973 3574 987 3578
rect 957 3557 961 3574
rect 983 3557 987 3574
rect 957 3527 961 3553
rect 974 3527 978 3553
rect 983 3527 987 3553
rect 991 3541 995 3582
rect 999 3569 1005 3573
rect 1011 3569 1028 3573
rect 999 3558 1003 3569
rect 1024 3559 1028 3569
rect 991 3537 1002 3541
rect 1009 3533 1013 3553
rect 991 3529 1013 3533
rect 974 3520 978 3523
rect 991 3520 995 3529
rect 1009 3527 1013 3529
rect 974 3516 995 3520
rect 1033 3542 1037 3553
rect 1033 3538 1036 3542
rect 1033 3527 1037 3538
rect 999 3519 1003 3522
rect 999 3516 1011 3519
rect 1024 3519 1028 3522
rect 1016 3516 1028 3519
rect 1001 3498 1004 3509
rect 898 3495 1004 3498
rect 194 3477 248 3481
rect 194 3442 197 3477
rect 207 3459 217 3463
rect 227 3463 264 3466
rect 269 3463 297 3466
rect 234 3460 238 3463
rect 252 3460 256 3463
rect 141 3438 197 3442
rect 276 3460 280 3463
rect 243 3443 247 3453
rect 286 3443 290 3455
rect 243 3439 278 3443
rect 286 3442 299 3443
rect 286 3439 318 3442
rect 142 3167 147 3438
rect 194 3434 197 3438
rect 233 3434 245 3435
rect 194 3431 245 3434
rect 252 3428 256 3439
rect 286 3429 290 3439
rect 295 3438 318 3439
rect 234 3419 238 3423
rect 276 3419 280 3422
rect 230 3416 289 3419
rect 315 3407 318 3438
rect 354 3440 357 3488
rect 757 3484 811 3488
rect 545 3476 591 3479
rect 597 3476 624 3479
rect 418 3469 456 3472
rect 550 3473 554 3476
rect 461 3469 483 3472
rect 606 3473 610 3476
rect 420 3466 424 3469
rect 438 3466 442 3469
rect 462 3466 466 3469
rect 429 3449 433 3459
rect 472 3449 476 3461
rect 540 3452 562 3455
rect 429 3445 464 3449
rect 472 3448 521 3449
rect 573 3448 577 3466
rect 616 3448 620 3468
rect 757 3453 760 3484
rect 790 3470 827 3473
rect 832 3470 860 3473
rect 797 3467 801 3470
rect 768 3462 778 3466
rect 815 3467 819 3470
rect 701 3448 760 3453
rect 472 3447 532 3448
rect 472 3445 552 3447
rect 417 3440 431 3441
rect 354 3437 431 3440
rect 438 3434 442 3445
rect 472 3435 476 3445
rect 518 3444 552 3445
rect 530 3443 552 3444
rect 560 3444 608 3448
rect 616 3444 624 3448
rect 420 3425 424 3429
rect 560 3434 564 3444
rect 416 3422 454 3425
rect 462 3425 466 3428
rect 616 3434 620 3444
rect 459 3422 477 3425
rect 550 3424 554 3428
rect 573 3424 577 3429
rect 545 3421 588 3424
rect 606 3424 610 3427
rect 594 3421 624 3424
rect 415 3353 422 3368
rect 701 3341 706 3448
rect 757 3441 760 3448
rect 839 3467 843 3470
rect 806 3450 810 3460
rect 849 3450 853 3462
rect 806 3446 841 3450
rect 849 3449 862 3450
rect 849 3446 881 3449
rect 796 3441 808 3442
rect 757 3438 808 3441
rect 815 3435 819 3446
rect 849 3436 853 3446
rect 858 3445 881 3446
rect 797 3426 801 3430
rect 839 3426 843 3429
rect 793 3423 852 3426
rect 878 3414 881 3445
rect 917 3447 920 3495
rect 1108 3483 1154 3486
rect 1160 3483 1187 3486
rect 981 3476 1019 3479
rect 1113 3480 1117 3483
rect 1024 3476 1046 3479
rect 1169 3480 1173 3483
rect 983 3473 987 3476
rect 1001 3473 1005 3476
rect 1025 3473 1029 3476
rect 992 3456 996 3466
rect 1035 3456 1039 3468
rect 1103 3459 1125 3462
rect 992 3452 1027 3456
rect 1035 3455 1084 3456
rect 1136 3455 1140 3473
rect 1179 3455 1183 3475
rect 1224 3455 1228 3609
rect 1335 3606 1341 3618
rect 1544 3614 1626 3619
rect 1619 3586 1626 3614
rect 1347 3567 1394 3571
rect 1347 3542 1351 3567
rect 1347 3512 1351 3538
rect 1356 3559 1371 3563
rect 1375 3559 1386 3563
rect 1356 3542 1360 3559
rect 1382 3542 1386 3559
rect 1356 3512 1360 3538
rect 1373 3512 1377 3538
rect 1382 3512 1386 3538
rect 1390 3526 1394 3567
rect 1398 3554 1415 3558
rect 1421 3554 1427 3558
rect 1398 3543 1402 3554
rect 1423 3544 1427 3554
rect 1390 3522 1401 3526
rect 1408 3518 1412 3538
rect 1390 3514 1412 3518
rect 1373 3505 1377 3508
rect 1390 3505 1394 3514
rect 1408 3512 1412 3514
rect 1373 3501 1394 3505
rect 1432 3527 1436 3538
rect 1432 3523 1435 3527
rect 1432 3512 1436 3523
rect 1398 3503 1401 3507
rect 1398 3500 1416 3503
rect 1424 3503 1427 3507
rect 1421 3500 1427 3503
rect 1384 3474 1387 3494
rect 1474 3484 1478 3574
rect 1524 3568 1571 3572
rect 1524 3543 1528 3568
rect 1524 3513 1528 3539
rect 1533 3560 1545 3564
rect 1549 3560 1563 3564
rect 1533 3543 1537 3560
rect 1559 3543 1563 3560
rect 1533 3513 1537 3539
rect 1550 3513 1554 3539
rect 1559 3513 1563 3539
rect 1567 3527 1571 3568
rect 1575 3555 1581 3559
rect 1587 3555 1604 3559
rect 1575 3544 1579 3555
rect 1600 3545 1604 3555
rect 1567 3523 1578 3527
rect 1585 3519 1589 3539
rect 1567 3515 1589 3519
rect 1550 3506 1554 3509
rect 1567 3506 1571 3515
rect 1585 3513 1589 3515
rect 1550 3502 1571 3506
rect 1609 3528 1613 3539
rect 1609 3524 1612 3528
rect 1609 3513 1613 3524
rect 1575 3505 1579 3508
rect 1575 3502 1587 3505
rect 1600 3505 1604 3508
rect 1592 3502 1604 3505
rect 1577 3484 1580 3495
rect 1474 3481 1580 3484
rect 1035 3454 1095 3455
rect 1035 3452 1115 3454
rect 980 3447 994 3448
rect 917 3444 994 3447
rect 1001 3441 1005 3452
rect 1035 3442 1039 3452
rect 1081 3451 1115 3452
rect 1093 3450 1115 3451
rect 1123 3451 1171 3455
rect 1179 3451 1228 3455
rect 1333 3470 1387 3474
rect 983 3432 987 3436
rect 1123 3441 1127 3451
rect 979 3429 1017 3432
rect 1025 3432 1029 3435
rect 1179 3441 1183 3451
rect 1022 3429 1040 3432
rect 1113 3431 1117 3435
rect 1136 3431 1140 3436
rect 1108 3428 1151 3431
rect 1169 3431 1173 3434
rect 1311 3431 1315 3432
rect 1333 3431 1336 3470
rect 1366 3456 1403 3459
rect 1408 3456 1436 3459
rect 1373 3453 1377 3456
rect 1345 3446 1353 3451
rect 1391 3453 1395 3456
rect 1415 3453 1419 3456
rect 1382 3436 1386 3446
rect 1425 3436 1429 3448
rect 1382 3432 1417 3436
rect 1425 3435 1438 3436
rect 1425 3432 1457 3435
rect 1157 3428 1187 3431
rect 1311 3427 1336 3431
rect 1372 3427 1384 3428
rect 902 3353 908 3373
rect 1218 3341 1223 3342
rect 700 3337 1223 3341
rect 174 3294 1079 3303
rect 174 3293 179 3294
rect 1075 3131 1079 3294
rect 1218 3146 1223 3337
rect 1311 3290 1315 3427
rect 1333 3424 1384 3427
rect 1391 3421 1395 3432
rect 1425 3422 1429 3432
rect 1434 3431 1457 3432
rect 1373 3412 1377 3416
rect 1415 3412 1419 3415
rect 1369 3409 1428 3412
rect 1454 3400 1457 3431
rect 1493 3433 1496 3481
rect 1684 3469 1730 3472
rect 1736 3469 1763 3472
rect 1557 3462 1595 3465
rect 1689 3466 1693 3469
rect 1600 3462 1622 3465
rect 1745 3466 1749 3469
rect 1559 3459 1563 3462
rect 1577 3459 1581 3462
rect 1601 3459 1605 3462
rect 1568 3442 1572 3452
rect 1611 3442 1615 3454
rect 1679 3445 1701 3448
rect 1568 3438 1603 3442
rect 1611 3441 1660 3442
rect 1712 3441 1716 3459
rect 1755 3441 1759 3461
rect 1783 3442 1789 3634
rect 1968 3598 2015 3602
rect 1968 3573 1972 3598
rect 1968 3543 1972 3569
rect 1977 3590 1992 3594
rect 1996 3590 2007 3594
rect 1977 3573 1981 3590
rect 2003 3573 2007 3590
rect 1977 3543 1981 3569
rect 1994 3543 1998 3569
rect 2003 3543 2007 3569
rect 2011 3557 2015 3598
rect 2019 3585 2036 3589
rect 2042 3585 2048 3589
rect 2019 3574 2023 3585
rect 2044 3575 2048 3585
rect 2011 3553 2022 3557
rect 2029 3549 2033 3569
rect 2011 3545 2033 3549
rect 1994 3536 1998 3539
rect 2011 3536 2015 3545
rect 2029 3543 2033 3545
rect 1994 3532 2015 3536
rect 2053 3558 2057 3569
rect 2053 3554 2056 3558
rect 2053 3543 2057 3554
rect 2019 3534 2022 3538
rect 2019 3531 2037 3534
rect 2045 3534 2048 3538
rect 2042 3531 2048 3534
rect 2005 3505 2008 3525
rect 2095 3515 2099 3605
rect 2145 3599 2192 3603
rect 2145 3574 2149 3599
rect 2145 3544 2149 3570
rect 2154 3591 2166 3595
rect 2170 3591 2184 3595
rect 2154 3574 2158 3591
rect 2180 3574 2184 3591
rect 2154 3544 2158 3570
rect 2171 3544 2175 3570
rect 2180 3544 2184 3570
rect 2188 3558 2192 3599
rect 2196 3586 2202 3590
rect 2208 3586 2225 3590
rect 2196 3575 2200 3586
rect 2221 3576 2225 3586
rect 2188 3554 2199 3558
rect 2206 3550 2210 3570
rect 2188 3546 2210 3550
rect 2171 3537 2175 3540
rect 2188 3537 2192 3546
rect 2206 3544 2210 3546
rect 2171 3533 2192 3537
rect 2230 3559 2234 3570
rect 2230 3555 2233 3559
rect 2264 3557 2414 3562
rect 2230 3544 2234 3555
rect 2196 3536 2200 3539
rect 2196 3533 2208 3536
rect 2221 3536 2225 3539
rect 2213 3533 2225 3536
rect 2198 3515 2201 3526
rect 2095 3512 2201 3515
rect 1939 3501 2008 3505
rect 1939 3469 1942 3501
rect 1955 3486 1964 3493
rect 1987 3487 2024 3490
rect 2029 3487 2057 3490
rect 1994 3484 1998 3487
rect 2012 3484 2016 3487
rect 1914 3464 1942 3469
rect 1762 3441 1789 3442
rect 1611 3440 1671 3441
rect 1611 3438 1691 3440
rect 1556 3433 1570 3434
rect 1493 3430 1570 3433
rect 1577 3427 1581 3438
rect 1611 3428 1615 3438
rect 1657 3437 1691 3438
rect 1669 3436 1691 3437
rect 1699 3437 1747 3441
rect 1755 3437 1789 3441
rect 1559 3418 1563 3422
rect 1699 3427 1703 3437
rect 1555 3415 1593 3418
rect 1601 3418 1605 3421
rect 1755 3427 1759 3437
rect 1598 3415 1616 3418
rect 1689 3417 1693 3421
rect 1712 3417 1716 3422
rect 1684 3414 1727 3417
rect 1745 3417 1749 3420
rect 1733 3414 1763 3417
rect 1557 3352 1563 3361
rect 1382 3290 1386 3291
rect 1311 3285 1386 3290
rect 1382 3170 1386 3285
rect 1552 3111 1557 3112
rect 1915 3111 1920 3464
rect 1939 3458 1942 3464
rect 2036 3484 2040 3487
rect 2003 3467 2007 3477
rect 2046 3467 2050 3479
rect 2003 3463 2038 3467
rect 2046 3466 2059 3467
rect 2046 3463 2078 3466
rect 1993 3458 2005 3459
rect 1939 3455 2005 3458
rect 2012 3452 2016 3463
rect 2046 3453 2050 3463
rect 2055 3462 2078 3463
rect 1994 3443 1998 3447
rect 2036 3443 2040 3446
rect 1990 3440 2049 3443
rect 2075 3431 2078 3462
rect 2114 3464 2117 3512
rect 2305 3500 2351 3503
rect 2357 3500 2384 3503
rect 2178 3493 2216 3496
rect 2310 3497 2314 3500
rect 2221 3493 2243 3496
rect 2366 3497 2370 3500
rect 2180 3490 2184 3493
rect 2198 3490 2202 3493
rect 2222 3490 2226 3493
rect 2189 3473 2193 3483
rect 2232 3473 2236 3485
rect 2300 3476 2322 3479
rect 2189 3469 2224 3473
rect 2232 3472 2281 3473
rect 2333 3472 2337 3490
rect 2376 3472 2380 3492
rect 2444 3472 2448 3670
rect 2232 3471 2292 3472
rect 2232 3469 2312 3471
rect 2177 3464 2191 3465
rect 2114 3461 2191 3464
rect 2198 3458 2202 3469
rect 2232 3459 2236 3469
rect 2278 3468 2312 3469
rect 2290 3467 2312 3468
rect 2320 3468 2368 3472
rect 2376 3468 2449 3472
rect 2180 3449 2184 3453
rect 2320 3458 2324 3468
rect 2176 3446 2214 3449
rect 2222 3449 2226 3452
rect 2376 3458 2380 3468
rect 2219 3446 2237 3449
rect 2310 3448 2314 3452
rect 2333 3448 2337 3453
rect 3380 3453 5023 3454
rect 2305 3445 2348 3448
rect 2366 3448 2370 3451
rect 2559 3448 5023 3453
rect 2354 3445 2384 3448
rect 2559 3447 3386 3448
rect 2086 3374 2093 3391
rect 1552 3106 1920 3111
rect 2255 3319 2260 3321
rect 2559 3319 2564 3447
rect 2255 3314 2566 3319
rect 2967 3316 2972 3421
rect 5015 3396 5021 3448
rect 4301 3370 5205 3376
rect 3162 3363 3168 3364
rect 3157 3357 3979 3363
rect 3162 3334 3168 3357
rect 3725 3339 3730 3340
rect 3161 3328 3238 3334
rect 316 3079 320 3081
rect 316 3076 1424 3079
rect 316 3044 320 3076
rect 382 3063 426 3066
rect 430 3063 458 3066
rect 395 3060 399 3063
rect 413 3060 417 3063
rect 437 3060 441 3063
rect 316 3040 397 3044
rect 404 3043 408 3053
rect 447 3043 451 3055
rect 230 2995 268 2998
rect 272 2995 305 2998
rect 237 2992 241 2995
rect 255 2992 259 2995
rect 279 2992 283 2995
rect 68 2972 239 2976
rect 246 2975 250 2985
rect 289 2975 293 2987
rect 68 2874 72 2972
rect 246 2971 281 2975
rect 289 2971 296 2975
rect 216 2963 248 2967
rect 173 2949 190 2952
rect 184 2942 205 2945
rect 190 2938 193 2942
rect 197 2925 201 2934
rect 216 2925 220 2963
rect 255 2960 259 2971
rect 289 2961 293 2971
rect 237 2951 241 2955
rect 279 2951 283 2954
rect 232 2948 295 2951
rect 300 2948 301 2951
rect 85 2921 186 2925
rect 197 2921 220 2925
rect 85 2902 89 2921
rect 197 2915 201 2921
rect 95 2911 131 2914
rect 100 2908 104 2911
rect 118 2908 122 2911
rect 135 2911 163 2914
rect 88 2897 89 2902
rect 85 2892 89 2897
rect 142 2908 146 2911
rect 190 2907 193 2911
rect 85 2888 102 2892
rect 109 2891 113 2901
rect 152 2891 156 2903
rect 174 2904 205 2907
rect 109 2887 144 2891
rect 152 2887 162 2891
rect 85 2879 111 2883
rect 85 2874 89 2879
rect 118 2876 122 2887
rect 68 2870 89 2874
rect 85 2842 89 2870
rect 152 2877 156 2887
rect 100 2864 104 2871
rect 142 2864 146 2870
rect 97 2861 157 2864
rect 174 2849 177 2904
rect 216 2895 220 2921
rect 227 2914 266 2917
rect 270 2914 297 2917
rect 236 2911 240 2914
rect 254 2911 258 2914
rect 278 2911 282 2914
rect 216 2891 238 2895
rect 245 2894 249 2904
rect 288 2894 292 2906
rect 316 2894 320 3040
rect 404 3039 439 3043
rect 447 3039 478 3043
rect 391 3031 406 3035
rect 413 3028 417 3039
rect 447 3029 451 3039
rect 500 3044 505 3076
rect 525 3063 569 3066
rect 573 3063 601 3066
rect 538 3060 542 3063
rect 556 3060 560 3063
rect 580 3060 584 3063
rect 500 3040 540 3044
rect 547 3043 551 3053
rect 590 3043 594 3055
rect 547 3039 582 3043
rect 590 3039 620 3043
rect 534 3031 549 3035
rect 395 3019 399 3023
rect 556 3028 560 3039
rect 437 3019 441 3022
rect 590 3029 594 3039
rect 663 3044 668 3076
rect 688 3063 732 3066
rect 736 3063 764 3066
rect 701 3060 705 3063
rect 719 3060 723 3063
rect 743 3060 747 3063
rect 663 3040 703 3044
rect 710 3043 714 3053
rect 753 3043 757 3055
rect 767 3043 780 3044
rect 710 3039 745 3043
rect 753 3039 780 3043
rect 819 3044 824 3076
rect 844 3063 888 3066
rect 892 3063 920 3066
rect 857 3060 861 3063
rect 875 3060 879 3063
rect 899 3060 903 3063
rect 819 3040 859 3044
rect 866 3043 870 3053
rect 909 3043 913 3055
rect 922 3043 931 3044
rect 866 3039 901 3043
rect 909 3039 931 3043
rect 956 3044 960 3076
rect 982 3063 1026 3066
rect 1030 3063 1058 3066
rect 995 3060 999 3063
rect 1013 3060 1017 3063
rect 1037 3060 1041 3063
rect 956 3040 997 3044
rect 1004 3043 1008 3053
rect 1047 3043 1051 3055
rect 1004 3039 1039 3043
rect 1047 3039 1074 3043
rect 1100 3044 1105 3076
rect 1125 3063 1169 3066
rect 1173 3063 1201 3066
rect 1138 3060 1142 3063
rect 1156 3060 1160 3063
rect 1180 3060 1184 3063
rect 1100 3040 1140 3044
rect 1147 3043 1151 3053
rect 1190 3043 1194 3055
rect 1147 3039 1182 3043
rect 1190 3039 1217 3043
rect 1263 3044 1268 3076
rect 1288 3063 1332 3066
rect 1336 3063 1364 3066
rect 1301 3060 1305 3063
rect 1319 3060 1323 3063
rect 1343 3060 1347 3063
rect 1263 3040 1303 3044
rect 1310 3043 1314 3053
rect 1353 3043 1357 3055
rect 1310 3039 1345 3043
rect 1353 3039 1380 3043
rect 697 3031 712 3035
rect 538 3019 542 3023
rect 719 3028 723 3039
rect 580 3019 584 3022
rect 753 3029 757 3039
rect 853 3031 868 3035
rect 701 3019 705 3023
rect 875 3028 879 3039
rect 743 3019 747 3022
rect 909 3029 913 3039
rect 991 3031 1006 3035
rect 857 3019 861 3023
rect 1013 3028 1017 3039
rect 899 3019 903 3022
rect 1047 3029 1051 3039
rect 1134 3031 1149 3035
rect 995 3019 999 3023
rect 1156 3028 1160 3039
rect 1037 3019 1041 3022
rect 1190 3029 1194 3039
rect 1297 3031 1312 3035
rect 1138 3019 1142 3023
rect 1319 3028 1323 3039
rect 1180 3019 1184 3022
rect 1353 3029 1357 3039
rect 1419 3044 1424 3076
rect 1444 3063 1488 3066
rect 1492 3063 1520 3066
rect 1457 3060 1461 3063
rect 1475 3060 1479 3063
rect 1499 3060 1503 3063
rect 1419 3040 1459 3044
rect 1466 3043 1470 3053
rect 1509 3043 1513 3055
rect 1552 3043 1557 3106
rect 1466 3039 1501 3043
rect 1509 3039 1557 3043
rect 1453 3031 1468 3035
rect 1301 3019 1305 3023
rect 1475 3028 1479 3039
rect 1343 3019 1347 3022
rect 1509 3029 1513 3039
rect 1457 3019 1461 3023
rect 1499 3019 1503 3022
rect 395 3016 455 3019
rect 538 3016 598 3019
rect 701 3016 761 3019
rect 857 3016 917 3019
rect 995 3016 1055 3019
rect 1138 3016 1198 3019
rect 1301 3016 1361 3019
rect 1457 3016 1517 3019
rect 426 3012 430 3016
rect 569 3012 573 3016
rect 732 3012 736 3016
rect 888 3012 892 3016
rect 1026 3012 1030 3016
rect 1169 3012 1173 3016
rect 1332 3012 1336 3016
rect 1488 3013 1492 3016
rect 1473 3012 1541 3013
rect 392 3008 1541 3012
rect 570 3007 659 3008
rect 729 3007 815 3008
rect 1170 3007 1259 3008
rect 1329 3007 1415 3008
rect 1488 3007 1491 3008
rect 1532 3007 1541 3008
rect 1552 3007 1554 3013
rect 2255 2991 2260 3314
rect 3232 3293 3238 3328
rect 3551 3319 3559 3339
rect 3723 3334 4123 3339
rect 3725 3328 3730 3334
rect 3725 3323 3795 3328
rect 3791 3298 3795 3323
rect 4301 3319 4307 3370
rect 4330 3334 4331 3339
rect 4340 3334 4546 3339
rect 4743 3338 4748 3348
rect 2965 3274 3012 3278
rect 2965 3249 2969 3274
rect 2965 3219 2969 3245
rect 2974 3266 2989 3270
rect 2993 3266 3004 3270
rect 2974 3249 2978 3266
rect 3000 3249 3004 3266
rect 2974 3219 2978 3245
rect 2991 3219 2995 3245
rect 3000 3219 3004 3245
rect 3008 3233 3012 3274
rect 3016 3261 3033 3265
rect 3039 3261 3045 3265
rect 3016 3250 3020 3261
rect 3041 3251 3045 3261
rect 3008 3229 3019 3233
rect 3026 3225 3030 3245
rect 3008 3221 3030 3225
rect 2991 3212 2995 3215
rect 3008 3212 3012 3221
rect 3026 3219 3030 3221
rect 2991 3208 3012 3212
rect 3050 3234 3054 3245
rect 3050 3230 3053 3234
rect 3050 3219 3054 3230
rect 3016 3210 3019 3214
rect 3016 3207 3034 3210
rect 3042 3210 3045 3214
rect 3039 3207 3045 3210
rect 3002 3181 3005 3201
rect 3092 3191 3096 3281
rect 3528 3281 3575 3285
rect 3142 3275 3189 3279
rect 3142 3250 3146 3275
rect 3142 3220 3146 3246
rect 3151 3267 3163 3271
rect 3167 3267 3181 3271
rect 3151 3250 3155 3267
rect 3177 3250 3181 3267
rect 3151 3220 3155 3246
rect 3168 3220 3172 3246
rect 3177 3220 3181 3246
rect 3185 3234 3189 3275
rect 3193 3262 3199 3266
rect 3205 3262 3222 3266
rect 3193 3251 3197 3262
rect 3218 3252 3222 3262
rect 3528 3256 3532 3281
rect 3185 3230 3196 3234
rect 3203 3226 3207 3246
rect 3185 3222 3207 3226
rect 3168 3213 3172 3216
rect 3185 3213 3189 3222
rect 3203 3220 3207 3222
rect 3168 3209 3189 3213
rect 3227 3235 3231 3246
rect 3227 3231 3230 3235
rect 3227 3220 3231 3231
rect 3528 3226 3532 3252
rect 3537 3273 3552 3277
rect 3556 3273 3567 3277
rect 3537 3256 3541 3273
rect 3563 3256 3567 3273
rect 3537 3226 3541 3252
rect 3554 3226 3558 3252
rect 3563 3226 3567 3252
rect 3571 3240 3575 3281
rect 3579 3268 3596 3272
rect 3602 3268 3608 3272
rect 3579 3257 3583 3268
rect 3604 3258 3608 3268
rect 3571 3236 3582 3240
rect 3589 3232 3593 3252
rect 3571 3228 3593 3232
rect 3193 3212 3197 3215
rect 3554 3219 3558 3222
rect 3571 3219 3575 3228
rect 3589 3226 3593 3228
rect 3554 3215 3575 3219
rect 3613 3241 3617 3252
rect 3613 3237 3616 3241
rect 3613 3226 3617 3237
rect 3579 3217 3582 3221
rect 3193 3209 3205 3212
rect 3218 3212 3222 3215
rect 3579 3214 3597 3217
rect 3605 3217 3608 3221
rect 3602 3214 3608 3217
rect 3210 3209 3222 3212
rect 3195 3191 3198 3202
rect 3092 3188 3198 3191
rect 3565 3188 3568 3208
rect 3655 3198 3659 3288
rect 3705 3282 3752 3286
rect 3705 3257 3709 3282
rect 3705 3227 3709 3253
rect 3714 3274 3726 3278
rect 3730 3274 3744 3278
rect 3714 3257 3718 3274
rect 3740 3257 3744 3274
rect 3714 3227 3718 3253
rect 3731 3227 3735 3253
rect 3740 3227 3744 3253
rect 3748 3241 3752 3282
rect 3756 3269 3762 3273
rect 3768 3269 3785 3273
rect 3756 3258 3760 3269
rect 3781 3259 3785 3269
rect 3748 3237 3759 3241
rect 3766 3233 3770 3253
rect 3748 3229 3770 3233
rect 3731 3220 3735 3223
rect 3748 3220 3752 3229
rect 3766 3227 3770 3229
rect 3731 3216 3752 3220
rect 3790 3242 3794 3253
rect 3790 3238 3793 3242
rect 3790 3227 3794 3238
rect 3756 3219 3760 3222
rect 3756 3216 3768 3219
rect 3781 3219 3785 3222
rect 3773 3216 3785 3219
rect 3758 3198 3761 3209
rect 3655 3195 3761 3198
rect 2951 3177 3005 3181
rect 2951 3142 2954 3177
rect 2964 3159 2974 3163
rect 2984 3163 3021 3166
rect 3026 3163 3054 3166
rect 2991 3160 2995 3163
rect 3009 3160 3013 3163
rect 2898 3138 2954 3142
rect 3033 3160 3037 3163
rect 3000 3143 3004 3153
rect 3043 3143 3047 3155
rect 3000 3139 3035 3143
rect 3043 3142 3056 3143
rect 3043 3139 3075 3142
rect 2379 2991 2381 2992
rect 1770 2990 1967 2991
rect 2176 2990 2381 2991
rect 1616 2989 1652 2990
rect 1659 2989 2381 2990
rect 1616 2987 2381 2989
rect 1616 2985 1784 2987
rect 1866 2986 2381 2987
rect 1616 2937 1620 2985
rect 1646 2984 1680 2985
rect 1635 2968 1696 2972
rect 1692 2964 1739 2968
rect 1692 2939 1696 2964
rect 245 2890 280 2894
rect 288 2890 320 2894
rect 337 2934 1621 2937
rect 337 2902 342 2934
rect 382 2921 426 2924
rect 430 2921 458 2924
rect 395 2918 399 2921
rect 413 2918 417 2921
rect 437 2918 441 2921
rect 337 2898 397 2902
rect 404 2901 408 2911
rect 447 2901 451 2913
rect 500 2902 505 2934
rect 525 2921 569 2924
rect 573 2921 601 2924
rect 538 2918 542 2921
rect 556 2918 560 2921
rect 580 2918 584 2921
rect 222 2882 247 2886
rect 184 2859 206 2862
rect 190 2855 193 2859
rect 197 2842 201 2851
rect 222 2842 226 2882
rect 254 2879 258 2890
rect 288 2880 292 2890
rect 236 2870 240 2874
rect 278 2870 282 2873
rect 234 2867 292 2870
rect 85 2838 186 2842
rect 197 2838 226 2842
rect 197 2833 201 2838
rect 190 2825 193 2829
rect 163 2819 166 2822
rect 185 2822 204 2825
rect 163 2738 167 2812
rect 215 2804 219 2838
rect 231 2823 270 2826
rect 274 2823 301 2826
rect 240 2820 244 2823
rect 258 2820 262 2823
rect 282 2820 286 2823
rect 215 2800 242 2804
rect 249 2803 253 2813
rect 292 2803 296 2815
rect 337 2803 342 2898
rect 404 2897 439 2901
rect 447 2897 467 2901
rect 391 2889 406 2893
rect 413 2886 417 2897
rect 447 2887 451 2897
rect 500 2898 540 2902
rect 547 2901 551 2911
rect 590 2901 594 2913
rect 602 2901 618 2902
rect 547 2897 582 2901
rect 590 2897 618 2901
rect 534 2889 549 2893
rect 395 2877 399 2881
rect 556 2886 560 2897
rect 437 2877 441 2880
rect 590 2887 594 2897
rect 663 2902 668 2934
rect 688 2921 732 2924
rect 736 2921 764 2924
rect 701 2918 705 2921
rect 719 2918 723 2921
rect 743 2918 747 2921
rect 663 2898 703 2902
rect 710 2901 714 2911
rect 753 2901 757 2913
rect 710 2897 745 2901
rect 753 2897 779 2901
rect 697 2889 712 2893
rect 538 2877 542 2881
rect 719 2886 723 2897
rect 580 2877 584 2880
rect 753 2887 757 2897
rect 819 2902 824 2934
rect 844 2921 888 2924
rect 892 2921 920 2924
rect 857 2918 861 2921
rect 875 2918 879 2921
rect 899 2918 903 2921
rect 819 2898 859 2902
rect 866 2901 870 2911
rect 909 2901 913 2913
rect 866 2897 901 2901
rect 909 2897 935 2901
rect 853 2889 868 2893
rect 701 2877 705 2881
rect 875 2886 879 2897
rect 743 2877 747 2880
rect 909 2887 913 2897
rect 956 2902 960 2934
rect 982 2921 1026 2924
rect 1030 2921 1058 2924
rect 995 2918 999 2921
rect 1013 2918 1017 2921
rect 1037 2918 1041 2921
rect 956 2898 997 2902
rect 1004 2901 1008 2911
rect 1047 2901 1051 2913
rect 1004 2897 1039 2901
rect 1047 2897 1074 2901
rect 991 2889 1006 2893
rect 857 2877 861 2881
rect 1013 2886 1017 2897
rect 899 2877 903 2880
rect 1047 2887 1051 2897
rect 1100 2902 1105 2934
rect 1125 2921 1169 2924
rect 1173 2921 1201 2924
rect 1138 2918 1142 2921
rect 1156 2918 1160 2921
rect 1180 2918 1184 2921
rect 1100 2898 1140 2902
rect 1147 2901 1151 2911
rect 1190 2901 1194 2913
rect 1147 2897 1182 2901
rect 1190 2897 1215 2901
rect 1263 2902 1268 2934
rect 1288 2921 1332 2924
rect 1336 2921 1364 2924
rect 1301 2918 1305 2921
rect 1319 2918 1323 2921
rect 1343 2918 1347 2921
rect 1263 2898 1303 2902
rect 1310 2901 1314 2911
rect 1353 2901 1357 2913
rect 1419 2902 1424 2934
rect 1444 2921 1488 2924
rect 1492 2921 1520 2924
rect 1589 2922 1624 2926
rect 1457 2918 1461 2921
rect 1475 2918 1479 2921
rect 1499 2918 1503 2921
rect 1310 2897 1345 2901
rect 1353 2897 1372 2901
rect 1134 2889 1149 2893
rect 995 2877 999 2881
rect 1156 2886 1160 2897
rect 1037 2877 1041 2880
rect 1190 2887 1194 2897
rect 1297 2889 1312 2893
rect 1138 2877 1142 2881
rect 1319 2886 1323 2897
rect 1180 2877 1184 2880
rect 1353 2887 1357 2897
rect 1419 2898 1459 2902
rect 1466 2901 1470 2911
rect 1509 2901 1513 2913
rect 1589 2901 1594 2922
rect 1692 2909 1696 2935
rect 1701 2956 1714 2960
rect 1720 2956 1731 2960
rect 1701 2939 1705 2956
rect 1727 2939 1731 2956
rect 1701 2909 1705 2935
rect 1718 2909 1722 2935
rect 1727 2909 1731 2935
rect 1735 2923 1739 2964
rect 1755 2955 1758 2976
rect 1772 2964 1779 2985
rect 1865 2971 1891 2974
rect 1887 2969 1891 2971
rect 1887 2965 1934 2969
rect 1743 2951 1772 2955
rect 1743 2940 1747 2951
rect 1768 2941 1772 2951
rect 1887 2940 1891 2965
rect 1735 2919 1746 2923
rect 1753 2915 1757 2935
rect 1735 2911 1757 2915
rect 1466 2897 1501 2901
rect 1509 2897 1594 2901
rect 1718 2902 1722 2905
rect 1735 2902 1739 2911
rect 1753 2909 1757 2911
rect 1718 2898 1739 2902
rect 1777 2924 1781 2935
rect 1777 2920 1780 2924
rect 1777 2909 1781 2920
rect 1743 2901 1747 2904
rect 1887 2910 1891 2936
rect 1896 2957 1906 2961
rect 1896 2940 1900 2957
rect 1912 2957 1926 2961
rect 1922 2940 1926 2957
rect 1896 2910 1900 2936
rect 1913 2910 1917 2936
rect 1922 2910 1926 2936
rect 1930 2924 1934 2965
rect 1950 2956 1953 2977
rect 1968 2965 1974 2986
rect 2079 2985 2194 2986
rect 2163 2981 2168 2982
rect 2072 2964 2147 2968
rect 1938 2952 1967 2956
rect 1938 2941 1942 2952
rect 1963 2942 1967 2952
rect 1930 2920 1941 2924
rect 1948 2916 1952 2936
rect 1930 2912 1952 2916
rect 1768 2901 1772 2904
rect 1743 2897 1772 2901
rect 1913 2903 1917 2906
rect 1930 2903 1934 2912
rect 1948 2910 1952 2912
rect 1913 2899 1934 2903
rect 1972 2925 1976 2936
rect 1972 2921 1975 2925
rect 1972 2910 1976 2921
rect 1938 2902 1942 2905
rect 2072 2907 2075 2964
rect 2100 2939 2104 2964
rect 2100 2909 2104 2935
rect 1963 2902 1967 2905
rect 1938 2898 1967 2902
rect 2109 2956 2121 2960
rect 2109 2939 2113 2956
rect 2128 2956 2139 2960
rect 2135 2939 2139 2956
rect 2109 2909 2113 2935
rect 2126 2909 2130 2935
rect 2135 2909 2139 2935
rect 2143 2923 2147 2964
rect 2163 2955 2166 2976
rect 2181 2967 2186 2985
rect 2284 2965 2348 2969
rect 2151 2951 2180 2955
rect 2151 2940 2155 2951
rect 2176 2941 2180 2951
rect 2301 2940 2305 2965
rect 2143 2919 2154 2923
rect 2161 2915 2165 2935
rect 2143 2911 2165 2915
rect 2126 2902 2130 2905
rect 2143 2902 2147 2911
rect 2161 2909 2165 2911
rect 2126 2898 2147 2902
rect 2185 2924 2189 2935
rect 2185 2920 2188 2924
rect 2185 2909 2189 2920
rect 2151 2901 2155 2904
rect 2301 2910 2305 2936
rect 2310 2957 2320 2961
rect 2326 2957 2340 2961
rect 2310 2940 2314 2957
rect 2336 2940 2340 2957
rect 2310 2910 2314 2936
rect 2327 2910 2331 2936
rect 2336 2910 2340 2936
rect 2344 2924 2348 2965
rect 2364 2956 2367 2977
rect 2352 2952 2381 2956
rect 2352 2941 2356 2952
rect 2377 2942 2381 2952
rect 2344 2920 2355 2924
rect 2362 2916 2366 2936
rect 2344 2912 2366 2916
rect 2176 2901 2180 2904
rect 1453 2889 1468 2893
rect 1301 2877 1305 2881
rect 1475 2886 1479 2897
rect 1343 2877 1347 2880
rect 1509 2887 1513 2897
rect 1457 2877 1461 2881
rect 1759 2883 1763 2897
rect 1954 2883 1958 2898
rect 2151 2897 2180 2901
rect 2327 2903 2331 2906
rect 2344 2903 2348 2912
rect 2362 2910 2366 2912
rect 2327 2899 2348 2903
rect 2386 2925 2390 2936
rect 2386 2921 2389 2925
rect 2386 2910 2390 2921
rect 2352 2902 2356 2905
rect 2377 2902 2381 2905
rect 2352 2898 2381 2902
rect 2167 2883 2171 2897
rect 2368 2883 2372 2898
rect 1759 2882 1958 2883
rect 2166 2882 2636 2883
rect 1499 2877 1503 2880
rect 1585 2879 2636 2882
rect 1585 2878 1872 2879
rect 2079 2878 2301 2879
rect 1585 2877 1592 2878
rect 2648 2879 2657 2883
rect 395 2874 455 2877
rect 538 2874 598 2877
rect 701 2874 761 2877
rect 857 2874 917 2877
rect 995 2874 1055 2877
rect 1138 2874 1198 2877
rect 1301 2874 1361 2877
rect 1457 2874 1592 2877
rect 426 2870 430 2874
rect 569 2870 573 2874
rect 732 2870 736 2874
rect 888 2870 892 2874
rect 1026 2870 1030 2874
rect 1169 2870 1173 2874
rect 1332 2870 1336 2874
rect 1488 2870 1492 2874
rect 392 2866 1492 2870
rect 570 2865 659 2866
rect 729 2865 815 2866
rect 1170 2865 1216 2866
rect 1231 2865 1259 2866
rect 1329 2865 1415 2866
rect 1380 2851 2071 2855
rect 249 2799 284 2803
rect 292 2799 343 2803
rect 2899 2800 2904 3138
rect 2951 3134 2954 3138
rect 2990 3134 3002 3135
rect 2951 3131 3002 3134
rect 3009 3128 3013 3139
rect 3043 3129 3047 3139
rect 3052 3138 3075 3139
rect 2991 3119 2995 3123
rect 3033 3119 3037 3122
rect 2987 3116 3046 3119
rect 3072 3107 3075 3138
rect 3111 3140 3114 3188
rect 3514 3184 3568 3188
rect 3302 3176 3348 3179
rect 3354 3176 3381 3179
rect 3175 3169 3213 3172
rect 3307 3173 3311 3176
rect 3218 3169 3240 3172
rect 3363 3173 3367 3176
rect 3177 3166 3181 3169
rect 3195 3166 3199 3169
rect 3219 3166 3223 3169
rect 3186 3149 3190 3159
rect 3229 3149 3233 3161
rect 3297 3152 3319 3155
rect 3186 3145 3221 3149
rect 3229 3148 3278 3149
rect 3330 3148 3334 3166
rect 3373 3148 3377 3168
rect 3514 3153 3517 3184
rect 3547 3170 3584 3173
rect 3589 3170 3617 3173
rect 3554 3167 3558 3170
rect 3525 3162 3535 3166
rect 3572 3167 3576 3170
rect 3458 3148 3517 3153
rect 3229 3147 3289 3148
rect 3229 3145 3309 3147
rect 3174 3140 3188 3141
rect 3111 3137 3188 3140
rect 3195 3134 3199 3145
rect 3229 3135 3233 3145
rect 3275 3144 3309 3145
rect 3287 3143 3309 3144
rect 3317 3144 3365 3148
rect 3373 3144 3381 3148
rect 3177 3125 3181 3129
rect 3317 3134 3321 3144
rect 3173 3122 3211 3125
rect 3219 3125 3223 3128
rect 3373 3134 3377 3144
rect 3216 3122 3234 3125
rect 3307 3124 3311 3128
rect 3330 3124 3334 3129
rect 3302 3121 3345 3124
rect 3363 3124 3367 3127
rect 3351 3121 3381 3124
rect 3172 3053 3179 3068
rect 2915 3036 2973 3041
rect 3458 2810 3463 3148
rect 3514 3141 3517 3148
rect 3596 3167 3600 3170
rect 3563 3150 3567 3160
rect 3606 3150 3610 3162
rect 3563 3146 3598 3150
rect 3606 3149 3619 3150
rect 3606 3146 3638 3149
rect 3553 3141 3565 3142
rect 3514 3138 3565 3141
rect 3572 3135 3576 3146
rect 3606 3136 3610 3146
rect 3615 3145 3638 3146
rect 3554 3126 3558 3130
rect 3596 3126 3600 3129
rect 3550 3123 3609 3126
rect 3635 3114 3638 3145
rect 3674 3147 3677 3195
rect 3865 3183 3911 3186
rect 3917 3183 3944 3186
rect 3738 3176 3776 3179
rect 3870 3180 3874 3183
rect 3781 3176 3803 3179
rect 3926 3180 3930 3183
rect 3740 3173 3744 3176
rect 3758 3173 3762 3176
rect 3782 3173 3786 3176
rect 3749 3156 3753 3166
rect 3792 3156 3796 3168
rect 3860 3159 3882 3162
rect 3749 3152 3784 3156
rect 3792 3155 3841 3156
rect 3893 3155 3897 3173
rect 3936 3155 3940 3175
rect 3981 3155 3985 3309
rect 4092 3306 4098 3318
rect 4301 3314 4383 3319
rect 4376 3286 4383 3314
rect 4104 3267 4151 3271
rect 4104 3242 4108 3267
rect 4104 3212 4108 3238
rect 4113 3259 4128 3263
rect 4132 3259 4143 3263
rect 4113 3242 4117 3259
rect 4139 3242 4143 3259
rect 4113 3212 4117 3238
rect 4130 3212 4134 3238
rect 4139 3212 4143 3238
rect 4147 3226 4151 3267
rect 4155 3254 4172 3258
rect 4178 3254 4184 3258
rect 4155 3243 4159 3254
rect 4180 3244 4184 3254
rect 4147 3222 4158 3226
rect 4165 3218 4169 3238
rect 4147 3214 4169 3218
rect 4130 3205 4134 3208
rect 4147 3205 4151 3214
rect 4165 3212 4169 3214
rect 4130 3201 4151 3205
rect 4189 3227 4193 3238
rect 4189 3223 4192 3227
rect 4189 3212 4193 3223
rect 4155 3203 4158 3207
rect 4155 3200 4173 3203
rect 4181 3203 4184 3207
rect 4178 3200 4184 3203
rect 4141 3174 4144 3194
rect 4231 3184 4235 3274
rect 4281 3268 4328 3272
rect 4281 3243 4285 3268
rect 4281 3213 4285 3239
rect 4290 3260 4302 3264
rect 4306 3260 4320 3264
rect 4290 3243 4294 3260
rect 4316 3243 4320 3260
rect 4290 3213 4294 3239
rect 4307 3213 4311 3239
rect 4316 3213 4320 3239
rect 4324 3227 4328 3268
rect 4332 3255 4338 3259
rect 4344 3255 4361 3259
rect 4332 3244 4336 3255
rect 4357 3245 4361 3255
rect 4324 3223 4335 3227
rect 4342 3219 4346 3239
rect 4324 3215 4346 3219
rect 4307 3206 4311 3209
rect 4324 3206 4328 3215
rect 4342 3213 4346 3215
rect 4307 3202 4328 3206
rect 4366 3228 4370 3239
rect 4366 3224 4369 3228
rect 4366 3213 4370 3224
rect 4332 3205 4336 3208
rect 4332 3202 4344 3205
rect 4357 3205 4361 3208
rect 4349 3202 4361 3205
rect 4334 3184 4337 3195
rect 4231 3181 4337 3184
rect 3792 3154 3852 3155
rect 3792 3152 3872 3154
rect 3737 3147 3751 3148
rect 3674 3144 3751 3147
rect 3758 3141 3762 3152
rect 3792 3142 3796 3152
rect 3838 3151 3872 3152
rect 3850 3150 3872 3151
rect 3880 3151 3928 3155
rect 3936 3151 3985 3155
rect 4090 3170 4144 3174
rect 3740 3132 3744 3136
rect 3880 3141 3884 3151
rect 3736 3129 3774 3132
rect 3782 3132 3786 3135
rect 3936 3141 3940 3151
rect 3779 3129 3797 3132
rect 3870 3131 3874 3135
rect 3893 3131 3897 3136
rect 3865 3128 3908 3131
rect 3926 3131 3930 3134
rect 4068 3131 4072 3132
rect 4090 3131 4093 3170
rect 4123 3156 4160 3159
rect 4165 3156 4193 3159
rect 4130 3153 4134 3156
rect 4102 3146 4110 3151
rect 4148 3153 4152 3156
rect 4172 3153 4176 3156
rect 4139 3136 4143 3146
rect 4182 3136 4186 3148
rect 4139 3132 4174 3136
rect 4182 3135 4195 3136
rect 4182 3132 4214 3135
rect 3914 3128 3944 3131
rect 4068 3127 4093 3131
rect 4129 3127 4141 3128
rect 3659 3053 3665 3073
rect 4068 3032 4072 3127
rect 4090 3124 4141 3127
rect 4148 3121 4152 3132
rect 4182 3122 4186 3132
rect 4191 3131 4214 3132
rect 4130 3112 4134 3116
rect 4172 3112 4176 3115
rect 4126 3109 4185 3112
rect 4211 3100 4214 3131
rect 4250 3133 4253 3181
rect 4441 3169 4487 3172
rect 4493 3169 4520 3172
rect 4314 3162 4352 3165
rect 4446 3166 4450 3169
rect 4357 3162 4379 3165
rect 4502 3166 4506 3169
rect 4316 3159 4320 3162
rect 4334 3159 4338 3162
rect 4358 3159 4362 3162
rect 4325 3142 4329 3152
rect 4368 3142 4372 3154
rect 4436 3145 4458 3148
rect 4325 3138 4360 3142
rect 4368 3141 4417 3142
rect 4469 3141 4473 3159
rect 4512 3141 4516 3161
rect 4540 3142 4546 3334
rect 4725 3298 4772 3302
rect 4725 3273 4729 3298
rect 4725 3243 4729 3269
rect 4734 3290 4749 3294
rect 4753 3290 4764 3294
rect 4734 3273 4738 3290
rect 4760 3273 4764 3290
rect 4734 3243 4738 3269
rect 4751 3243 4755 3269
rect 4760 3243 4764 3269
rect 4768 3257 4772 3298
rect 4776 3285 4793 3289
rect 4799 3285 4805 3289
rect 4776 3274 4780 3285
rect 4801 3275 4805 3285
rect 4768 3253 4779 3257
rect 4786 3249 4790 3269
rect 4768 3245 4790 3249
rect 4751 3236 4755 3239
rect 4768 3236 4772 3245
rect 4786 3243 4790 3245
rect 4751 3232 4772 3236
rect 4810 3258 4814 3269
rect 4810 3254 4813 3258
rect 4810 3243 4814 3254
rect 4776 3234 4779 3238
rect 4776 3231 4794 3234
rect 4802 3234 4805 3238
rect 4799 3231 4805 3234
rect 4762 3205 4765 3225
rect 4852 3215 4856 3305
rect 4902 3299 4949 3303
rect 4902 3274 4906 3299
rect 4902 3244 4906 3270
rect 4911 3291 4923 3295
rect 4927 3291 4941 3295
rect 4911 3274 4915 3291
rect 4937 3274 4941 3291
rect 4911 3244 4915 3270
rect 4928 3244 4932 3270
rect 4937 3244 4941 3270
rect 4945 3258 4949 3299
rect 4953 3286 4959 3290
rect 4965 3286 4982 3290
rect 4953 3275 4957 3286
rect 4978 3276 4982 3286
rect 4945 3254 4956 3258
rect 4963 3250 4967 3270
rect 4945 3246 4967 3250
rect 4928 3237 4932 3240
rect 4945 3237 4949 3246
rect 4963 3244 4967 3246
rect 4928 3233 4949 3237
rect 4987 3259 4991 3270
rect 4987 3255 4990 3259
rect 4987 3244 4991 3255
rect 4953 3236 4957 3239
rect 4953 3233 4965 3236
rect 4978 3236 4982 3239
rect 4970 3233 4982 3236
rect 4955 3215 4958 3226
rect 4852 3212 4958 3215
rect 4696 3201 4765 3205
rect 4696 3169 4699 3201
rect 4712 3186 4721 3193
rect 4744 3187 4781 3190
rect 4786 3187 4814 3190
rect 4751 3184 4755 3187
rect 4769 3184 4773 3187
rect 4671 3164 4699 3169
rect 4519 3141 4546 3142
rect 4368 3140 4428 3141
rect 4368 3138 4448 3140
rect 4313 3133 4327 3134
rect 4250 3130 4327 3133
rect 4334 3127 4338 3138
rect 4368 3128 4372 3138
rect 4414 3137 4448 3138
rect 4426 3136 4448 3137
rect 4456 3137 4504 3141
rect 4512 3137 4546 3141
rect 4316 3118 4320 3122
rect 4456 3127 4460 3137
rect 4312 3115 4350 3118
rect 4358 3118 4362 3121
rect 4512 3127 4516 3137
rect 4355 3115 4373 3118
rect 4446 3117 4450 3121
rect 4469 3117 4473 3122
rect 4441 3114 4484 3117
rect 4502 3117 4506 3120
rect 4490 3114 4520 3117
rect 4314 3052 4320 3061
rect 4068 2825 4073 3032
rect 4672 2841 4677 3164
rect 4696 3158 4699 3164
rect 4793 3184 4797 3187
rect 4760 3167 4764 3177
rect 4803 3167 4807 3179
rect 4760 3163 4795 3167
rect 4803 3166 4816 3167
rect 4803 3163 4835 3166
rect 4750 3158 4762 3159
rect 4696 3155 4762 3158
rect 4769 3152 4773 3163
rect 4803 3153 4807 3163
rect 4812 3162 4835 3163
rect 4751 3143 4755 3147
rect 4793 3143 4797 3146
rect 4747 3140 4806 3143
rect 4832 3131 4835 3162
rect 4871 3164 4874 3212
rect 5062 3200 5108 3203
rect 5114 3200 5141 3203
rect 4935 3193 4973 3196
rect 5067 3197 5071 3200
rect 4978 3193 5000 3196
rect 5123 3197 5127 3200
rect 4937 3190 4941 3193
rect 4955 3190 4959 3193
rect 4979 3190 4983 3193
rect 4946 3173 4950 3183
rect 4989 3173 4993 3185
rect 5057 3176 5079 3179
rect 4946 3169 4981 3173
rect 4989 3172 5038 3173
rect 5090 3172 5094 3190
rect 5133 3172 5137 3192
rect 5201 3172 5205 3370
rect 4989 3171 5049 3172
rect 4989 3169 5069 3171
rect 4934 3164 4948 3165
rect 4871 3161 4948 3164
rect 4955 3158 4959 3169
rect 4989 3159 4993 3169
rect 5035 3168 5069 3169
rect 5047 3167 5069 3168
rect 5077 3168 5125 3172
rect 5133 3168 5206 3172
rect 4937 3149 4941 3153
rect 5077 3158 5081 3168
rect 4933 3146 4971 3149
rect 4979 3149 4983 3152
rect 5133 3158 5137 3168
rect 4976 3146 4994 3149
rect 5067 3148 5071 3152
rect 5090 3148 5094 3153
rect 5062 3145 5105 3148
rect 5123 3148 5127 3151
rect 5111 3145 5141 3148
rect 4843 3074 4850 3091
rect 236 2791 251 2795
rect 258 2788 262 2799
rect 292 2789 296 2799
rect 240 2779 244 2783
rect 347 2785 1813 2788
rect 282 2779 286 2782
rect 238 2776 296 2779
rect 347 2760 351 2785
rect 382 2772 426 2775
rect 430 2772 458 2775
rect 395 2769 399 2772
rect 413 2769 417 2772
rect 291 2754 351 2760
rect 347 2753 351 2754
rect 437 2769 441 2772
rect 347 2749 397 2753
rect 404 2752 408 2762
rect 447 2752 451 2764
rect 500 2753 505 2785
rect 525 2772 569 2775
rect 573 2772 601 2775
rect 538 2769 542 2772
rect 556 2769 560 2772
rect 580 2769 584 2772
rect 404 2748 439 2752
rect 447 2748 476 2752
rect 500 2749 540 2753
rect 547 2752 551 2762
rect 590 2752 594 2764
rect 663 2753 668 2785
rect 688 2772 732 2775
rect 736 2772 764 2775
rect 701 2769 705 2772
rect 719 2769 723 2772
rect 743 2769 747 2772
rect 547 2748 582 2752
rect 590 2748 614 2752
rect 663 2749 703 2753
rect 710 2752 714 2762
rect 753 2752 757 2764
rect 819 2753 824 2785
rect 844 2772 888 2775
rect 892 2772 920 2775
rect 857 2769 861 2772
rect 875 2769 879 2772
rect 899 2769 903 2772
rect 710 2748 745 2752
rect 753 2748 783 2752
rect 819 2749 859 2753
rect 866 2752 870 2762
rect 909 2752 913 2764
rect 956 2753 960 2785
rect 982 2772 1026 2775
rect 1030 2772 1058 2775
rect 995 2769 999 2772
rect 1013 2769 1017 2772
rect 1037 2769 1041 2772
rect 866 2748 901 2752
rect 909 2748 937 2752
rect 956 2749 997 2753
rect 1004 2752 1008 2762
rect 1047 2752 1051 2764
rect 1100 2753 1105 2785
rect 1125 2772 1169 2775
rect 1173 2772 1201 2775
rect 1138 2769 1142 2772
rect 1156 2769 1160 2772
rect 1180 2769 1184 2772
rect 1004 2748 1039 2752
rect 1047 2748 1082 2752
rect 391 2740 406 2744
rect 162 2646 166 2738
rect 413 2737 417 2748
rect 447 2738 451 2748
rect 534 2740 549 2744
rect 395 2728 399 2732
rect 556 2737 560 2748
rect 437 2728 441 2731
rect 590 2738 594 2748
rect 697 2740 712 2744
rect 538 2728 542 2732
rect 719 2737 723 2748
rect 580 2728 584 2731
rect 753 2738 757 2748
rect 853 2740 868 2744
rect 701 2728 705 2732
rect 875 2737 879 2748
rect 743 2728 747 2731
rect 909 2738 913 2748
rect 991 2740 1006 2744
rect 857 2728 861 2732
rect 1013 2737 1017 2748
rect 899 2728 903 2731
rect 1047 2738 1051 2748
rect 1100 2749 1140 2753
rect 1147 2752 1151 2762
rect 1190 2752 1194 2764
rect 1263 2753 1268 2785
rect 1288 2772 1332 2775
rect 1336 2772 1364 2775
rect 1301 2769 1305 2772
rect 1319 2769 1323 2772
rect 1343 2769 1347 2772
rect 1147 2748 1182 2752
rect 1190 2748 1227 2752
rect 1263 2749 1303 2753
rect 1310 2752 1314 2762
rect 1353 2752 1357 2764
rect 1419 2753 1424 2785
rect 1444 2772 1488 2775
rect 1492 2772 1520 2775
rect 1457 2769 1461 2772
rect 1475 2769 1479 2772
rect 1499 2769 1503 2772
rect 1310 2748 1345 2752
rect 1353 2748 1365 2752
rect 1134 2740 1149 2744
rect 995 2728 999 2732
rect 1156 2737 1160 2748
rect 1037 2728 1041 2731
rect 1190 2738 1194 2748
rect 1297 2740 1312 2744
rect 1138 2728 1142 2732
rect 1319 2737 1323 2748
rect 1180 2728 1184 2731
rect 1353 2738 1357 2748
rect 1419 2749 1459 2753
rect 1466 2752 1470 2762
rect 1509 2752 1513 2764
rect 1809 2766 1812 2785
rect 2281 2778 2287 2785
rect 2281 2774 2967 2778
rect 2281 2766 2287 2774
rect 1809 2761 2288 2766
rect 2324 2756 2488 2759
rect 1466 2748 1501 2752
rect 1509 2748 1520 2752
rect 1453 2740 1468 2744
rect 1301 2728 1305 2732
rect 1475 2737 1479 2748
rect 1343 2728 1347 2731
rect 1509 2738 1513 2748
rect 1457 2728 1461 2732
rect 1499 2728 1503 2731
rect 395 2725 455 2728
rect 538 2725 598 2728
rect 701 2725 761 2728
rect 857 2725 917 2728
rect 995 2725 1055 2728
rect 1138 2725 1198 2728
rect 1301 2725 1361 2728
rect 1457 2725 1517 2728
rect 426 2721 430 2725
rect 569 2721 573 2725
rect 732 2721 736 2725
rect 888 2721 892 2725
rect 1026 2721 1030 2725
rect 1169 2721 1173 2725
rect 1332 2721 1336 2725
rect 1488 2721 1492 2725
rect 392 2717 2081 2721
rect 570 2716 659 2717
rect 729 2716 815 2717
rect 1170 2716 1259 2717
rect 1329 2716 1415 2717
rect 347 2660 1424 2663
rect 162 2635 167 2646
rect 347 2635 351 2660
rect 382 2647 426 2650
rect 430 2647 458 2650
rect 395 2644 399 2647
rect 413 2644 417 2647
rect 162 2629 351 2635
rect 347 2628 351 2629
rect 437 2644 441 2647
rect 347 2624 397 2628
rect 404 2627 408 2637
rect 447 2627 451 2639
rect 404 2623 439 2627
rect 447 2623 468 2627
rect 500 2628 505 2660
rect 525 2647 569 2650
rect 573 2647 601 2650
rect 538 2644 542 2647
rect 556 2644 560 2647
rect 580 2644 584 2647
rect 500 2624 540 2628
rect 547 2627 551 2637
rect 590 2627 594 2639
rect 663 2628 668 2660
rect 688 2647 732 2650
rect 736 2647 764 2650
rect 701 2644 705 2647
rect 719 2644 723 2647
rect 743 2644 747 2647
rect 547 2623 582 2627
rect 590 2623 612 2627
rect 391 2615 406 2619
rect 413 2612 417 2623
rect 447 2613 451 2623
rect 534 2615 549 2619
rect 395 2603 399 2607
rect 556 2612 560 2623
rect 437 2603 441 2606
rect 590 2613 594 2623
rect 663 2624 703 2628
rect 710 2627 714 2637
rect 753 2627 757 2639
rect 710 2623 745 2627
rect 753 2623 778 2627
rect 697 2615 712 2619
rect 538 2603 542 2607
rect 719 2612 723 2623
rect 580 2603 584 2606
rect 753 2613 757 2623
rect 819 2628 824 2660
rect 844 2647 888 2650
rect 892 2647 920 2650
rect 857 2644 861 2647
rect 875 2644 879 2647
rect 899 2644 903 2647
rect 819 2624 859 2628
rect 866 2627 870 2637
rect 909 2627 913 2639
rect 956 2628 960 2660
rect 982 2647 1026 2650
rect 1030 2647 1058 2650
rect 995 2644 999 2647
rect 1013 2644 1017 2647
rect 1037 2644 1041 2647
rect 866 2623 901 2627
rect 909 2623 922 2627
rect 853 2615 868 2619
rect 701 2603 705 2607
rect 875 2612 879 2623
rect 743 2603 747 2606
rect 909 2613 913 2623
rect 956 2624 997 2628
rect 1004 2627 1008 2637
rect 1047 2627 1051 2639
rect 1004 2623 1039 2627
rect 1047 2623 1067 2627
rect 991 2615 1006 2619
rect 857 2603 861 2607
rect 1013 2612 1017 2623
rect 899 2603 903 2606
rect 1047 2613 1051 2623
rect 1100 2628 1105 2660
rect 1125 2647 1169 2650
rect 1173 2647 1201 2650
rect 1138 2644 1142 2647
rect 1156 2644 1160 2647
rect 1180 2644 1184 2647
rect 1100 2624 1140 2628
rect 1147 2627 1151 2637
rect 1190 2627 1194 2639
rect 1147 2623 1182 2627
rect 1190 2623 1219 2627
rect 1134 2615 1149 2619
rect 995 2603 999 2607
rect 1156 2612 1160 2623
rect 1037 2603 1041 2606
rect 1190 2613 1194 2623
rect 1263 2628 1268 2660
rect 1288 2647 1332 2650
rect 1336 2647 1364 2650
rect 1301 2644 1305 2647
rect 1319 2644 1323 2647
rect 1343 2644 1347 2647
rect 1263 2624 1303 2628
rect 1310 2627 1314 2637
rect 1353 2627 1357 2639
rect 1310 2623 1345 2627
rect 1353 2623 1376 2627
rect 1297 2615 1312 2619
rect 1138 2603 1142 2607
rect 1319 2612 1323 2623
rect 1180 2603 1184 2606
rect 1353 2613 1357 2623
rect 1419 2628 1424 2660
rect 2073 2659 2077 2717
rect 2112 2697 2123 2701
rect 2128 2698 2164 2701
rect 2128 2697 2137 2698
rect 2118 2692 2121 2697
rect 2324 2701 2327 2756
rect 2360 2746 2364 2756
rect 2390 2746 2394 2756
rect 2420 2746 2424 2756
rect 2445 2746 2449 2756
rect 2373 2726 2377 2742
rect 2405 2726 2409 2742
rect 2435 2726 2439 2742
rect 2461 2726 2465 2742
rect 2373 2722 2452 2726
rect 2461 2722 2467 2726
rect 2435 2711 2439 2722
rect 2461 2717 2465 2722
rect 2172 2698 2327 2701
rect 2360 2701 2364 2707
rect 2445 2701 2449 2707
rect 2485 2707 2488 2756
rect 2485 2704 2874 2707
rect 2360 2698 2476 2701
rect 2126 2676 2129 2688
rect 2360 2686 2364 2698
rect 2161 2682 2364 2686
rect 2126 2672 2131 2676
rect 2126 2668 2129 2672
rect 2119 2659 2122 2664
rect 2161 2659 2164 2682
rect 2383 2681 2387 2684
rect 2398 2681 2402 2684
rect 2413 2681 2417 2684
rect 2427 2681 2431 2684
rect 2073 2656 2131 2659
rect 2073 2655 2121 2656
rect 2136 2656 2164 2659
rect 1444 2647 1488 2650
rect 1492 2647 1520 2650
rect 1457 2644 1461 2647
rect 1475 2644 1479 2647
rect 1499 2644 1503 2647
rect 1419 2624 1459 2628
rect 1466 2627 1470 2637
rect 1509 2627 1513 2639
rect 2114 2631 2122 2635
rect 2127 2631 2139 2635
rect 1466 2623 1501 2627
rect 1509 2623 1559 2627
rect 1453 2615 1468 2619
rect 1301 2603 1305 2607
rect 1475 2612 1479 2623
rect 1343 2603 1347 2606
rect 1509 2613 1513 2623
rect 1521 2622 1536 2623
rect 1457 2603 1461 2607
rect 1499 2603 1503 2606
rect 395 2600 455 2603
rect 538 2600 598 2603
rect 701 2600 761 2603
rect 857 2600 917 2603
rect 995 2600 1055 2603
rect 1138 2600 1198 2603
rect 1301 2600 1361 2603
rect 1457 2600 1517 2603
rect 239 2592 316 2596
rect 260 2237 267 2592
rect 326 2592 327 2596
rect 426 2596 430 2600
rect 569 2596 573 2600
rect 732 2596 736 2600
rect 888 2596 892 2600
rect 1026 2596 1030 2600
rect 1169 2596 1173 2600
rect 1332 2596 1336 2600
rect 1488 2596 1492 2600
rect 392 2592 1492 2596
rect 570 2591 659 2592
rect 729 2591 815 2592
rect 1170 2591 1259 2592
rect 1329 2591 1415 2592
rect 738 2452 1066 2461
rect 738 2269 742 2452
rect 882 2413 1221 2420
rect 764 2288 808 2291
rect 812 2288 840 2291
rect 777 2285 781 2288
rect 795 2285 799 2288
rect 819 2285 823 2288
rect 738 2265 779 2269
rect 786 2268 790 2278
rect 829 2268 833 2280
rect 882 2269 887 2413
rect 1045 2395 1050 2398
rect 1044 2390 1376 2395
rect 907 2288 951 2291
rect 955 2288 983 2291
rect 920 2285 924 2288
rect 938 2285 942 2288
rect 962 2285 966 2288
rect 786 2264 821 2268
rect 829 2264 846 2268
rect 882 2265 922 2269
rect 929 2268 933 2278
rect 972 2268 976 2280
rect 1045 2269 1050 2390
rect 1246 2389 1376 2390
rect 1554 2367 1559 2623
rect 2120 2626 2123 2631
rect 2128 2610 2131 2622
rect 2128 2606 2141 2610
rect 2128 2602 2131 2606
rect 2121 2593 2124 2598
rect 2473 2597 2476 2698
rect 2485 2659 2488 2704
rect 2810 2696 2814 2704
rect 2870 2696 2874 2704
rect 2862 2677 2866 2692
rect 2883 2681 2887 2692
rect 2883 2677 2892 2681
rect 2823 2673 2876 2677
rect 2823 2669 2827 2673
rect 2849 2669 2853 2673
rect 2883 2669 2887 2677
rect 2485 2656 2606 2659
rect 2491 2646 2495 2656
rect 2524 2646 2528 2656
rect 2553 2646 2557 2656
rect 2562 2646 2566 2656
rect 2506 2626 2511 2642
rect 2539 2626 2543 2642
rect 2578 2626 2582 2642
rect 2506 2622 2569 2626
rect 2578 2622 2584 2626
rect 2553 2611 2557 2622
rect 2578 2617 2582 2622
rect 2603 2621 2606 2656
rect 2810 2657 2814 2662
rect 2836 2657 2840 2662
rect 2862 2657 2866 2665
rect 2870 2657 2874 2665
rect 2810 2654 2874 2657
rect 2603 2618 2736 2621
rect 2491 2597 2495 2607
rect 2562 2597 2566 2607
rect 2629 2608 2633 2618
rect 2662 2608 2666 2618
rect 2688 2608 2692 2618
rect 2473 2594 2603 2597
rect 2120 2590 2131 2593
rect 2117 2564 2122 2568
rect 2127 2564 2142 2568
rect 2534 2571 2538 2584
rect 2402 2568 2538 2571
rect 2123 2559 2126 2564
rect 2544 2564 2548 2583
rect 2417 2561 2548 2564
rect 2600 2559 2603 2594
rect 2644 2588 2649 2604
rect 2679 2588 2683 2604
rect 2704 2588 2708 2604
rect 2644 2584 2695 2588
rect 2704 2584 2710 2588
rect 2679 2573 2683 2584
rect 2704 2579 2708 2584
rect 2733 2578 2736 2618
rect 2733 2574 2825 2578
rect 2629 2559 2633 2569
rect 2688 2559 2692 2569
rect 2758 2568 2762 2574
rect 2600 2556 2726 2559
rect 2131 2543 2134 2555
rect 2193 2546 2637 2550
rect 2193 2543 2197 2546
rect 2131 2539 2197 2543
rect 2131 2535 2134 2539
rect 2672 2537 2676 2545
rect 2403 2534 2676 2537
rect 2723 2531 2726 2556
rect 2769 2548 2773 2565
rect 2779 2568 2783 2574
rect 2806 2569 2809 2574
rect 2790 2548 2794 2565
rect 2814 2553 2817 2565
rect 2797 2549 2802 2553
rect 2814 2549 2818 2553
rect 2797 2548 2800 2549
rect 2769 2544 2800 2548
rect 2814 2545 2817 2549
rect 2758 2531 2762 2537
rect 2790 2538 2794 2544
rect 2807 2531 2810 2541
rect 2867 2531 2870 2654
rect 2124 2526 2127 2531
rect 2723 2528 2870 2531
rect 2123 2523 2131 2526
rect 2117 2497 2122 2501
rect 2127 2497 2142 2501
rect 2123 2492 2126 2497
rect 2131 2476 2134 2488
rect 2131 2472 2574 2476
rect 2131 2468 2134 2472
rect 2124 2459 2127 2464
rect 2123 2456 2131 2459
rect 2104 2392 2122 2396
rect 2041 2374 2081 2378
rect 1201 2363 1560 2367
rect 1070 2288 1114 2291
rect 1118 2288 1146 2291
rect 1083 2285 1087 2288
rect 1101 2285 1105 2288
rect 1125 2285 1129 2288
rect 929 2264 964 2268
rect 972 2264 989 2268
rect 1045 2265 1085 2269
rect 1092 2268 1096 2278
rect 1135 2268 1139 2280
rect 1201 2269 1206 2363
rect 1545 2362 1560 2363
rect 2041 2350 2045 2374
rect 2041 2333 2045 2346
rect 2028 2330 2045 2333
rect 2041 2319 2045 2330
rect 2050 2367 2069 2371
rect 2050 2350 2054 2367
rect 2069 2350 2073 2366
rect 2050 2319 2054 2346
rect 2060 2319 2064 2346
rect 2069 2319 2073 2346
rect 2077 2334 2081 2374
rect 2104 2366 2108 2392
rect 2127 2392 2160 2396
rect 2141 2387 2144 2392
rect 2149 2371 2152 2383
rect 2135 2367 2137 2371
rect 2149 2367 2259 2371
rect 2085 2362 2108 2366
rect 2149 2363 2152 2367
rect 2085 2350 2089 2362
rect 2104 2350 2108 2362
rect 2142 2354 2145 2359
rect 2130 2351 2145 2354
rect 2077 2330 2087 2334
rect 2094 2326 2098 2346
rect 2077 2322 2098 2326
rect 2060 2312 2064 2315
rect 2077 2312 2081 2322
rect 2094 2319 2098 2322
rect 2113 2334 2117 2346
rect 2113 2330 2116 2334
rect 2113 2319 2117 2330
rect 2060 2308 2081 2312
rect 2085 2312 2089 2315
rect 2104 2312 2108 2315
rect 2130 2313 2135 2351
rect 2130 2312 2131 2313
rect 2085 2308 2131 2312
rect 1946 2299 2010 2303
rect 2027 2301 2065 2304
rect 1226 2288 1270 2291
rect 2007 2291 2010 2299
rect 2027 2291 2030 2301
rect 1274 2288 1302 2291
rect 1973 2288 2030 2291
rect 1239 2285 1243 2288
rect 1257 2285 1261 2288
rect 1281 2285 1285 2288
rect 1092 2264 1127 2268
rect 1135 2264 1152 2268
rect 1201 2265 1241 2269
rect 1248 2268 1252 2278
rect 1291 2268 1295 2280
rect 1248 2264 1283 2268
rect 1291 2264 1308 2268
rect 773 2256 788 2260
rect 795 2253 799 2264
rect 829 2254 833 2264
rect 916 2256 931 2260
rect 777 2244 781 2248
rect 938 2253 942 2264
rect 819 2244 823 2247
rect 972 2254 976 2264
rect 1079 2256 1094 2260
rect 920 2244 924 2248
rect 1101 2253 1105 2264
rect 962 2244 966 2247
rect 1135 2254 1139 2264
rect 1235 2256 1250 2260
rect 1083 2244 1087 2248
rect 1257 2253 1261 2264
rect 1125 2244 1129 2247
rect 1291 2254 1295 2264
rect 1239 2244 1243 2248
rect 1281 2244 1285 2247
rect 777 2241 837 2244
rect 920 2241 980 2244
rect 1083 2241 1143 2244
rect 1239 2241 1299 2244
rect 808 2237 812 2241
rect 951 2237 955 2241
rect 1114 2237 1118 2241
rect 1270 2237 1274 2241
rect 260 2233 1274 2237
rect 952 2232 1041 2233
rect 1111 2232 1197 2233
rect 1884 2133 1943 2138
rect 1845 1980 1942 1984
rect 1951 1980 1953 1984
rect 1973 1544 1976 2288
rect 2106 2231 2122 2235
rect 2043 2213 2083 2217
rect 2043 2189 2047 2213
rect 2043 2172 2047 2185
rect 2030 2169 2047 2172
rect 2043 2158 2047 2169
rect 2052 2206 2071 2210
rect 2052 2189 2056 2206
rect 2071 2189 2075 2205
rect 2052 2158 2056 2185
rect 2062 2158 2066 2185
rect 2071 2158 2075 2185
rect 2079 2173 2083 2213
rect 2106 2205 2110 2231
rect 2127 2231 2157 2235
rect 2143 2226 2146 2231
rect 2151 2210 2154 2222
rect 2137 2206 2139 2210
rect 2151 2208 2221 2210
rect 2087 2201 2110 2205
rect 2151 2205 2222 2208
rect 2151 2202 2154 2205
rect 2087 2189 2091 2201
rect 2106 2189 2110 2201
rect 2144 2193 2147 2198
rect 2079 2169 2089 2173
rect 2096 2165 2100 2185
rect 2079 2161 2100 2165
rect 2062 2151 2066 2154
rect 2079 2151 2083 2161
rect 2096 2158 2100 2161
rect 2115 2173 2119 2185
rect 2137 2190 2147 2193
rect 2115 2169 2118 2173
rect 2115 2158 2119 2169
rect 2062 2147 2083 2151
rect 2087 2151 2091 2154
rect 2106 2151 2110 2154
rect 2132 2151 2137 2188
rect 2087 2147 2137 2151
rect 2029 2140 2067 2143
rect 2029 2133 2032 2140
rect 2213 2139 2222 2205
rect 2250 2159 2259 2367
rect 2652 2260 2656 2524
rect 2784 2512 2788 2519
rect 2962 2435 2967 2774
rect 2962 2292 2966 2435
rect 2304 2257 2656 2260
rect 2735 2182 2874 2185
rect 2738 2172 2742 2182
rect 2771 2172 2775 2182
rect 2800 2172 2804 2182
rect 2809 2172 2813 2182
rect 2871 2176 2874 2182
rect 2871 2173 2964 2176
rect 2250 2154 2397 2159
rect 2402 2154 2696 2159
rect 2251 2153 2696 2154
rect 1991 2130 2007 2133
rect 1991 1687 1994 2130
rect 2014 2130 2032 2133
rect 2213 2134 2412 2139
rect 2417 2134 2675 2139
rect 2213 2132 2675 2134
rect 2213 2131 2222 2132
rect 2672 2110 2675 2132
rect 2693 2117 2696 2153
rect 2753 2152 2758 2168
rect 2786 2152 2790 2168
rect 2825 2152 2829 2168
rect 2901 2170 2905 2173
rect 2921 2170 2925 2173
rect 2943 2170 2947 2173
rect 2912 2153 2916 2163
rect 2953 2153 2957 2165
rect 2753 2148 2816 2152
rect 2825 2148 2904 2152
rect 2800 2137 2804 2148
rect 2825 2143 2829 2148
rect 2912 2149 2945 2153
rect 2953 2149 2961 2153
rect 2920 2138 2924 2149
rect 2738 2123 2742 2133
rect 2809 2128 2813 2133
rect 2953 2139 2957 2149
rect 2901 2129 2905 2133
rect 2943 2129 2947 2132
rect 2893 2128 2961 2129
rect 2809 2126 2961 2128
rect 2809 2125 2896 2126
rect 2809 2123 2813 2125
rect 2738 2120 2808 2123
rect 2693 2114 2720 2117
rect 2672 2107 2720 2110
rect 2574 2099 2720 2102
rect 2047 2091 2058 2095
rect 2105 2077 2122 2081
rect 2042 2059 2082 2063
rect 2042 2035 2046 2059
rect 2042 2018 2046 2031
rect 2029 2015 2046 2018
rect 2042 2004 2046 2015
rect 2051 2052 2070 2056
rect 2051 2035 2055 2052
rect 2070 2035 2074 2051
rect 2051 2004 2055 2031
rect 2061 2004 2065 2031
rect 2070 2004 2074 2031
rect 2078 2019 2082 2059
rect 2105 2051 2109 2077
rect 2127 2077 2161 2081
rect 2142 2072 2145 2077
rect 2150 2056 2153 2068
rect 2136 2052 2138 2056
rect 2150 2052 2426 2056
rect 2574 2056 2577 2099
rect 2431 2052 2577 2056
rect 2646 2090 2720 2093
rect 2086 2047 2109 2051
rect 2150 2048 2153 2052
rect 2086 2035 2090 2047
rect 2105 2035 2109 2047
rect 2143 2039 2146 2044
rect 2078 2015 2088 2019
rect 2095 2011 2099 2031
rect 2078 2007 2099 2011
rect 2061 1997 2065 2000
rect 2078 1997 2082 2007
rect 2095 2004 2099 2007
rect 2114 2019 2118 2031
rect 2136 2036 2146 2039
rect 2114 2015 2117 2019
rect 2114 2004 2118 2015
rect 2061 1993 2082 1997
rect 2086 1997 2090 2000
rect 2105 1997 2109 2000
rect 2131 1997 2136 2034
rect 2086 1993 2136 1997
rect 2028 1986 2066 1989
rect 2028 1978 2031 1986
rect 2002 1975 2017 1978
rect 2002 1751 2005 1975
rect 2023 1975 2031 1978
rect 2105 1929 2122 1933
rect 2042 1911 2082 1915
rect 2042 1887 2046 1911
rect 2042 1870 2046 1883
rect 2029 1867 2046 1870
rect 2042 1856 2046 1867
rect 2051 1904 2070 1908
rect 2051 1887 2055 1904
rect 2070 1887 2074 1903
rect 2051 1856 2055 1883
rect 2061 1856 2065 1883
rect 2070 1856 2074 1883
rect 2078 1871 2082 1911
rect 2105 1903 2109 1929
rect 2127 1929 2161 1933
rect 2142 1924 2145 1929
rect 2150 1908 2153 1920
rect 2646 1908 2652 2090
rect 2136 1904 2138 1908
rect 2150 1904 2652 1908
rect 2742 1924 2865 1927
rect 2086 1899 2109 1903
rect 2150 1900 2153 1904
rect 2086 1887 2090 1899
rect 2105 1887 2109 1899
rect 2143 1891 2146 1896
rect 2078 1867 2088 1871
rect 2095 1863 2099 1883
rect 2078 1859 2099 1863
rect 2061 1849 2065 1852
rect 2078 1849 2082 1859
rect 2095 1856 2099 1859
rect 2114 1871 2118 1883
rect 2136 1888 2146 1891
rect 2114 1867 2117 1871
rect 2114 1856 2118 1867
rect 2061 1845 2082 1849
rect 2086 1849 2090 1852
rect 2105 1849 2109 1852
rect 2131 1849 2136 1886
rect 2742 1870 2745 1924
rect 2801 1916 2805 1924
rect 2861 1916 2865 1924
rect 2853 1897 2857 1912
rect 2874 1901 2878 1912
rect 2874 1897 2883 1901
rect 2814 1893 2867 1897
rect 2814 1889 2818 1893
rect 2840 1889 2844 1893
rect 2874 1889 2878 1897
rect 2801 1877 2805 1882
rect 2827 1877 2831 1882
rect 2853 1877 2857 1885
rect 2861 1877 2865 1885
rect 2801 1874 2865 1877
rect 2571 1867 2745 1870
rect 2575 1857 2579 1867
rect 2605 1857 2609 1867
rect 2635 1857 2639 1867
rect 2660 1857 2664 1867
rect 2086 1845 2136 1849
rect 2028 1838 2066 1841
rect 2028 1824 2031 1838
rect 2588 1837 2592 1853
rect 2620 1837 2624 1853
rect 2650 1837 2654 1853
rect 2676 1837 2680 1853
rect 2588 1833 2667 1837
rect 2676 1833 2682 1837
rect 2034 1821 2570 1824
rect 2650 1822 2654 1833
rect 2676 1828 2680 1833
rect 2112 1802 2122 1806
rect 2127 1802 2137 1806
rect 2118 1797 2121 1802
rect 2126 1781 2129 1793
rect 2537 1786 2540 1807
rect 2565 1791 2570 1821
rect 2575 1812 2579 1818
rect 2660 1812 2664 1818
rect 2814 1812 2817 1874
rect 2835 1859 2839 1865
rect 2575 1809 2817 1812
rect 2598 1791 2602 1794
rect 2565 1788 2602 1791
rect 2440 1783 2540 1786
rect 2082 1777 2101 1781
rect 2126 1777 2185 1781
rect 2126 1773 2129 1777
rect 2443 1773 2447 1783
rect 2476 1773 2480 1783
rect 2505 1773 2509 1783
rect 2514 1773 2518 1783
rect 2119 1764 2122 1769
rect 2118 1761 2131 1764
rect 2458 1753 2463 1769
rect 2491 1753 2495 1769
rect 2530 1753 2534 1769
rect 2002 1747 2425 1751
rect 2458 1749 2521 1753
rect 2530 1749 2536 1753
rect 2114 1736 2122 1740
rect 2127 1736 2139 1740
rect 2120 1731 2123 1736
rect 2128 1715 2131 1727
rect 2082 1711 2101 1715
rect 2128 1711 2142 1715
rect 2128 1707 2131 1711
rect 2299 1708 2383 1711
rect 2121 1698 2124 1703
rect 2302 1698 2306 1708
rect 2335 1698 2339 1708
rect 2361 1698 2365 1708
rect 2421 1707 2425 1747
rect 2505 1738 2509 1749
rect 2530 1744 2534 1749
rect 2443 1724 2447 1734
rect 2514 1724 2518 1734
rect 2605 1724 2608 1809
rect 2613 1786 2617 1794
rect 2443 1721 2608 1724
rect 2466 1707 2470 1711
rect 2421 1704 2470 1707
rect 2476 1699 2480 1721
rect 2486 1706 2490 1712
rect 2496 1706 2500 1712
rect 2120 1695 2131 1698
rect 1991 1684 2290 1687
rect 2117 1669 2122 1673
rect 2127 1669 2142 1673
rect 2123 1664 2126 1669
rect 2131 1648 2134 1660
rect 2074 1644 2101 1648
rect 2131 1644 2136 1648
rect 2131 1640 2134 1644
rect 2124 1631 2127 1636
rect 2123 1628 2131 1631
rect 2186 1630 2270 1634
rect 2117 1602 2122 1606
rect 2186 1606 2189 1630
rect 2207 1624 2211 1630
rect 2127 1602 2189 1606
rect 2218 1604 2222 1621
rect 2228 1624 2232 1630
rect 2255 1625 2258 1630
rect 2287 1630 2290 1684
rect 2317 1678 2322 1694
rect 2352 1678 2356 1694
rect 2377 1678 2381 1694
rect 2431 1696 2480 1699
rect 2317 1674 2368 1678
rect 2377 1674 2384 1678
rect 2352 1663 2356 1674
rect 2377 1669 2381 1674
rect 2302 1649 2306 1659
rect 2361 1649 2365 1659
rect 2431 1649 2434 1696
rect 2471 1685 2474 1687
rect 2628 1685 2632 1795
rect 2642 1787 2646 1795
rect 2471 1682 2632 1685
rect 2302 1646 2434 1649
rect 2325 1630 2329 1636
rect 2287 1627 2329 1630
rect 2239 1604 2243 1621
rect 2263 1609 2266 1621
rect 2246 1605 2251 1609
rect 2263 1605 2267 1609
rect 2246 1604 2249 1605
rect 2123 1597 2126 1602
rect 2218 1600 2249 1604
rect 2263 1601 2266 1605
rect 2131 1581 2134 1593
rect 2207 1586 2211 1593
rect 2239 1594 2243 1600
rect 2256 1586 2259 1597
rect 2336 1586 2339 1646
rect 2345 1631 2349 1635
rect 2207 1583 2339 1586
rect 2053 1577 2101 1581
rect 2131 1577 2137 1581
rect 2131 1573 2134 1577
rect 2124 1564 2127 1569
rect 2222 1564 2225 1583
rect 2123 1561 2131 1564
rect 2136 1561 2225 1564
rect 2233 1544 2237 1573
rect 1973 1541 2237 1544
<< m2contact >>
rect 1222 3655 1229 3664
rect 209 3604 221 3616
rect 1366 3632 1377 3642
rect 794 3608 803 3619
rect 1574 3631 1583 3642
rect 1222 3609 1229 3618
rect 276 3561 282 3567
rect 277 3506 282 3511
rect 442 3562 448 3568
rect 839 3568 845 3574
rect 448 3508 453 3513
rect 840 3513 845 3518
rect 1005 3569 1011 3575
rect 1011 3515 1016 3520
rect 200 3458 207 3464
rect 264 3463 269 3468
rect 289 3415 295 3420
rect 591 3476 597 3482
rect 413 3469 418 3474
rect 456 3469 461 3474
rect 827 3470 832 3475
rect 763 3462 768 3467
rect 454 3420 459 3426
rect 588 3420 594 3425
rect 415 3368 423 3377
rect 852 3422 858 3427
rect 1154 3483 1160 3489
rect 976 3476 981 3481
rect 1019 3476 1024 3481
rect 1335 3598 1343 3606
rect 1415 3554 1421 3560
rect 1416 3499 1421 3504
rect 1581 3555 1587 3561
rect 1587 3501 1592 3506
rect 1017 3427 1022 3433
rect 1151 3427 1157 3432
rect 1403 3456 1408 3461
rect 1339 3446 1345 3452
rect 902 3373 910 3381
rect 165 3293 174 3304
rect 139 3157 149 3167
rect 1428 3408 1434 3413
rect 1730 3469 1736 3475
rect 1552 3462 1557 3467
rect 1595 3462 1600 3467
rect 1985 3629 1993 3638
rect 2036 3585 2042 3591
rect 2037 3530 2042 3535
rect 2202 3586 2208 3592
rect 2414 3556 2420 3564
rect 2208 3532 2213 3537
rect 1946 3486 1955 3496
rect 2024 3487 2029 3492
rect 1593 3413 1598 3419
rect 1727 3413 1733 3418
rect 1557 3361 1565 3369
rect 1380 3161 1387 3170
rect 1215 3136 1224 3146
rect 1074 3120 1083 3131
rect 2049 3439 2055 3444
rect 2351 3500 2357 3506
rect 2173 3493 2178 3498
rect 2216 3493 2221 3498
rect 2214 3444 2219 3450
rect 2348 3444 2354 3449
rect 2086 3391 2096 3398
rect 3979 3355 3986 3364
rect 296 2971 301 2977
rect 295 2948 300 2953
rect 83 2897 88 2902
rect 162 2886 168 2893
rect 385 3030 391 3036
rect 478 3037 488 3047
rect 528 3030 534 3036
rect 620 3038 630 3048
rect 780 3039 785 3045
rect 931 3039 937 3046
rect 1074 3039 1081 3046
rect 1217 3039 1226 3049
rect 691 3030 697 3036
rect 847 3030 853 3036
rect 985 3030 991 3036
rect 1128 3030 1134 3036
rect 1291 3030 1297 3036
rect 1380 3038 1387 3047
rect 1447 3030 1453 3036
rect 386 3007 392 3013
rect 2966 3304 2978 3316
rect 4123 3332 4134 3342
rect 3551 3308 3560 3319
rect 4331 3331 4340 3342
rect 3979 3309 3986 3318
rect 3033 3261 3039 3267
rect 3034 3206 3039 3211
rect 3199 3262 3205 3268
rect 3596 3268 3602 3274
rect 3205 3208 3210 3213
rect 3597 3213 3602 3218
rect 3762 3269 3768 3275
rect 3768 3215 3773 3220
rect 2957 3158 2964 3164
rect 3021 3163 3026 3168
rect 1628 2967 1635 2974
rect 292 2867 297 2872
rect 163 2812 169 2819
rect 385 2888 391 2894
rect 467 2896 474 2902
rect 528 2888 534 2894
rect 618 2896 626 2903
rect 691 2888 697 2894
rect 779 2896 787 2903
rect 847 2888 853 2894
rect 935 2895 942 2903
rect 985 2888 991 2894
rect 1074 2895 1084 2904
rect 1215 2897 1222 2903
rect 1128 2888 1134 2894
rect 1291 2888 1297 2894
rect 1372 2896 1380 2902
rect 1714 2956 1720 2961
rect 1857 2968 1865 2975
rect 1906 2956 1912 2962
rect 2121 2955 2128 2961
rect 2320 2957 2326 2962
rect 1447 2888 1453 2894
rect 386 2865 392 2871
rect 1372 2850 1380 2856
rect 3046 3115 3052 3120
rect 3348 3176 3354 3182
rect 3170 3169 3175 3174
rect 3213 3169 3218 3174
rect 3584 3170 3589 3175
rect 3520 3162 3525 3167
rect 3211 3120 3216 3126
rect 3345 3120 3351 3125
rect 3172 3068 3180 3077
rect 2908 3035 2915 3041
rect 2973 3035 2981 3043
rect 3609 3122 3615 3127
rect 3911 3183 3917 3189
rect 3733 3176 3738 3181
rect 3776 3176 3781 3181
rect 4092 3298 4100 3306
rect 4172 3254 4178 3260
rect 4173 3199 4178 3204
rect 4338 3255 4344 3261
rect 4344 3201 4349 3206
rect 3774 3127 3779 3133
rect 3908 3127 3914 3132
rect 4160 3156 4165 3161
rect 4096 3146 4102 3152
rect 3659 3073 3667 3081
rect 4185 3108 4191 3113
rect 4487 3169 4493 3175
rect 4309 3162 4314 3167
rect 4352 3162 4357 3167
rect 4742 3329 4750 3338
rect 4793 3285 4799 3291
rect 4794 3230 4799 3235
rect 4959 3286 4965 3292
rect 4965 3232 4970 3237
rect 4703 3186 4712 3196
rect 4781 3187 4786 3192
rect 4350 3113 4355 3119
rect 4484 3113 4490 3118
rect 4314 3061 4322 3069
rect 4806 3139 4812 3144
rect 5108 3200 5114 3206
rect 4930 3193 4935 3198
rect 4973 3193 4978 3198
rect 4971 3144 4976 3150
rect 5105 3144 5111 3149
rect 4843 3091 4853 3098
rect 4669 2830 4681 2841
rect 4066 2815 4077 2825
rect 3458 2802 3467 2810
rect 228 2790 236 2797
rect 2897 2793 2907 2800
rect 296 2776 301 2781
rect 282 2754 291 2762
rect 476 2748 482 2753
rect 614 2748 620 2753
rect 783 2748 788 2753
rect 937 2748 944 2753
rect 385 2739 391 2745
rect 528 2739 534 2745
rect 691 2739 697 2745
rect 847 2739 853 2745
rect 985 2739 991 2745
rect 1082 2747 1087 2753
rect 1227 2748 1233 2753
rect 1128 2739 1134 2745
rect 1291 2739 1297 2745
rect 1365 2747 1372 2753
rect 1520 2748 1527 2753
rect 1447 2739 1453 2745
rect 386 2716 392 2722
rect 468 2623 474 2629
rect 385 2614 391 2620
rect 528 2614 534 2620
rect 612 2622 619 2628
rect 691 2614 697 2620
rect 778 2622 788 2630
rect 847 2614 853 2620
rect 922 2621 928 2628
rect 985 2614 991 2620
rect 1067 2622 1074 2629
rect 1128 2614 1134 2620
rect 1219 2621 1230 2629
rect 1291 2614 1297 2620
rect 1376 2620 1386 2631
rect 2382 2676 2387 2681
rect 2397 2676 2402 2681
rect 2412 2676 2417 2681
rect 2426 2676 2431 2681
rect 1447 2614 1453 2620
rect 316 2591 326 2599
rect 386 2591 392 2597
rect 1066 2450 1078 2461
rect 1221 2412 1233 2424
rect 1376 2387 1386 2398
rect 2397 2567 2402 2572
rect 2412 2560 2417 2565
rect 2398 2533 2403 2538
rect 2023 2328 2028 2333
rect 2069 2366 2074 2371
rect 2130 2367 2135 2372
rect 767 2255 773 2261
rect 910 2255 916 2261
rect 1073 2255 1079 2261
rect 1229 2255 1235 2261
rect 2025 2167 2030 2172
rect 2071 2205 2076 2210
rect 2132 2206 2137 2211
rect 2299 2255 2304 2260
rect 2397 2154 2402 2159
rect 2412 2134 2417 2139
rect 2042 2090 2047 2095
rect 2024 2013 2029 2018
rect 2070 2051 2075 2056
rect 2131 2052 2136 2057
rect 2426 2052 2431 2057
rect 2024 1865 2029 1870
rect 2070 1903 2075 1908
rect 2131 1904 2136 1909
rect 2566 1865 2571 1870
rect 2536 1807 2541 1812
rect 2077 1777 2082 1782
rect 2077 1710 2082 1715
rect 2294 1706 2299 1711
rect 2612 1781 2617 1786
rect 2485 1701 2490 1706
rect 2495 1701 2500 1706
rect 2069 1643 2074 1648
rect 2270 1629 2275 1634
rect 2469 1687 2474 1692
rect 2641 1782 2646 1787
rect 2345 1626 2350 1631
rect 2048 1576 2053 1581
<< metal2 >>
rect 182 3606 209 3611
rect 183 3587 188 3606
rect 745 3613 794 3618
rect 221 3606 619 3611
rect 183 3487 186 3587
rect 277 3567 281 3606
rect 400 3605 438 3606
rect 443 3568 447 3606
rect 516 3583 523 3606
rect 183 3484 269 3487
rect 264 3468 269 3484
rect 278 3484 282 3506
rect 448 3495 451 3508
rect 374 3492 451 3495
rect 278 3480 330 3484
rect 165 3463 171 3464
rect 164 3459 200 3463
rect 165 3304 171 3459
rect 284 3416 289 3419
rect 289 3373 293 3415
rect 327 3373 330 3480
rect 374 3373 378 3492
rect 517 3482 523 3583
rect 413 3479 523 3482
rect 591 3482 596 3606
rect 746 3594 751 3613
rect 1224 3618 1228 3655
rect 1377 3634 1574 3639
rect 1942 3630 1985 3635
rect 803 3613 1182 3618
rect 746 3494 749 3594
rect 840 3574 844 3613
rect 1006 3575 1010 3613
rect 1079 3590 1086 3613
rect 746 3491 832 3494
rect 413 3478 451 3479
rect 413 3474 416 3478
rect 456 3474 460 3479
rect 827 3475 832 3491
rect 841 3491 845 3513
rect 1011 3502 1014 3515
rect 937 3499 1014 3502
rect 841 3487 893 3491
rect 662 3462 763 3466
rect 456 3413 459 3420
rect 456 3409 480 3413
rect 187 3368 415 3373
rect 475 3373 480 3409
rect 588 3373 592 3420
rect 423 3368 621 3373
rect 327 3367 330 3368
rect 662 3283 667 3462
rect 847 3423 852 3426
rect 852 3380 856 3422
rect 890 3380 893 3487
rect 750 3375 902 3380
rect 890 3374 893 3375
rect 937 3380 941 3499
rect 1080 3489 1086 3590
rect 976 3486 1086 3489
rect 1154 3489 1159 3613
rect 1943 3611 1948 3630
rect 1993 3630 2379 3635
rect 1224 3607 1228 3609
rect 1321 3599 1335 3604
rect 1322 3580 1327 3599
rect 1343 3599 1758 3604
rect 976 3485 1014 3486
rect 976 3481 979 3485
rect 1019 3481 1023 3486
rect 1322 3480 1325 3580
rect 1416 3560 1420 3599
rect 1537 3598 1564 3599
rect 1582 3561 1586 3599
rect 1655 3576 1662 3599
rect 1322 3477 1408 3480
rect 1403 3461 1408 3477
rect 1417 3477 1421 3499
rect 1587 3488 1590 3501
rect 1513 3485 1590 3488
rect 1417 3473 1469 3477
rect 1291 3446 1339 3451
rect 1019 3420 1022 3427
rect 1019 3416 1043 3420
rect 1038 3380 1043 3416
rect 1151 3380 1155 3427
rect 910 3375 1184 3380
rect 621 3279 667 3283
rect 149 3158 483 3165
rect 480 3047 483 3158
rect 621 3048 625 3279
rect 780 3209 784 3211
rect 1292 3209 1296 3446
rect 1423 3409 1428 3412
rect 1428 3366 1432 3408
rect 1466 3366 1469 3473
rect 1513 3366 1517 3485
rect 1656 3475 1662 3576
rect 1552 3472 1662 3475
rect 1730 3475 1735 3599
rect 1943 3511 1946 3611
rect 2037 3591 2041 3630
rect 2203 3592 2207 3630
rect 2276 3607 2283 3630
rect 1943 3508 2029 3511
rect 1801 3493 1808 3494
rect 1801 3486 1946 3493
rect 2024 3492 2029 3508
rect 2038 3508 2042 3530
rect 2208 3519 2211 3532
rect 2134 3516 2211 3519
rect 2038 3504 2090 3508
rect 2085 3503 2090 3504
rect 1552 3471 1590 3472
rect 1552 3467 1555 3471
rect 1595 3467 1599 3472
rect 1595 3406 1598 3413
rect 1595 3402 1619 3406
rect 1326 3361 1557 3366
rect 1614 3366 1619 3402
rect 1727 3366 1731 3413
rect 1565 3361 1760 3366
rect 1466 3360 1469 3361
rect 779 3204 1296 3209
rect 780 3045 784 3204
rect 931 3188 935 3190
rect 1801 3188 1808 3486
rect 2044 3440 2049 3443
rect 2049 3397 2053 3439
rect 2087 3398 2090 3503
rect 1947 3392 2086 3397
rect 2134 3397 2138 3516
rect 2277 3506 2283 3607
rect 2173 3503 2283 3506
rect 2351 3506 2356 3630
rect 2173 3502 2211 3503
rect 2173 3498 2176 3502
rect 2216 3498 2220 3503
rect 2216 3437 2219 3444
rect 2216 3433 2240 3437
rect 2235 3397 2240 3433
rect 2348 3420 2352 3444
rect 2415 3420 2419 3556
rect 2348 3416 2422 3420
rect 2348 3397 2352 3416
rect 2096 3392 2381 3397
rect 2939 3306 2966 3311
rect 931 3183 1808 3188
rect 2940 3287 2945 3306
rect 3502 3313 3551 3318
rect 2978 3306 3376 3311
rect 2940 3187 2943 3287
rect 3034 3267 3038 3306
rect 3157 3305 3195 3306
rect 3200 3268 3204 3306
rect 3273 3283 3280 3306
rect 2940 3184 3026 3187
rect 931 3046 935 3183
rect 3021 3168 3026 3184
rect 3035 3184 3039 3206
rect 3205 3195 3208 3208
rect 3131 3192 3208 3195
rect 3035 3180 3087 3184
rect 2922 3163 2928 3164
rect 1075 3046 1079 3120
rect 1218 3049 1223 3136
rect 1382 3047 1386 3161
rect 2921 3159 2957 3163
rect 2922 3049 2928 3159
rect 3041 3116 3046 3119
rect 3046 3073 3050 3115
rect 3084 3073 3087 3180
rect 3131 3073 3135 3192
rect 3274 3182 3280 3283
rect 3170 3179 3280 3182
rect 3348 3182 3353 3306
rect 3503 3294 3508 3313
rect 3981 3318 3985 3355
rect 4134 3334 4331 3339
rect 4699 3330 4742 3335
rect 3560 3313 3939 3318
rect 3503 3194 3506 3294
rect 3597 3274 3601 3313
rect 3763 3275 3767 3313
rect 3836 3290 3843 3313
rect 3503 3191 3589 3194
rect 3170 3178 3208 3179
rect 3170 3174 3173 3178
rect 3213 3174 3217 3179
rect 3584 3175 3589 3191
rect 3598 3191 3602 3213
rect 3768 3202 3771 3215
rect 3694 3199 3771 3202
rect 3598 3187 3650 3191
rect 3419 3162 3520 3166
rect 3213 3113 3216 3120
rect 3213 3109 3237 3113
rect 2944 3068 3172 3073
rect 3232 3073 3237 3109
rect 3345 3073 3349 3120
rect 3180 3068 3378 3073
rect 3084 3067 3087 3068
rect 2216 3046 2928 3049
rect 2216 3037 2220 3046
rect 371 3031 385 3035
rect 391 3031 392 3035
rect 514 3031 528 3035
rect 534 3031 535 3035
rect 677 3031 691 3035
rect 697 3031 698 3035
rect 833 3031 847 3035
rect 853 3031 854 3035
rect 971 3031 985 3035
rect 991 3031 992 3035
rect 1114 3031 1128 3035
rect 1134 3031 1135 3035
rect 1277 3031 1291 3035
rect 1297 3031 1298 3035
rect 1433 3031 1447 3035
rect 1453 3031 1454 3035
rect 1714 3034 2220 3037
rect 2233 3036 2908 3041
rect 44 3013 49 3014
rect 44 3008 300 3013
rect 44 2760 49 3008
rect 296 2977 300 3008
rect 328 3008 386 3011
rect 328 2951 332 3008
rect 1590 2967 1628 2972
rect 1590 2955 1595 2967
rect 1714 2961 1718 3034
rect 2233 3025 2239 3036
rect 3419 3041 3424 3162
rect 3604 3123 3609 3126
rect 3609 3080 3613 3122
rect 3647 3080 3650 3187
rect 3507 3075 3659 3080
rect 3647 3074 3650 3075
rect 3694 3080 3698 3199
rect 3837 3189 3843 3290
rect 3733 3186 3843 3189
rect 3911 3189 3916 3313
rect 4700 3311 4705 3330
rect 4750 3330 5136 3335
rect 3981 3307 3985 3309
rect 4078 3299 4092 3304
rect 4079 3280 4084 3299
rect 4100 3299 4515 3304
rect 3733 3185 3771 3186
rect 3733 3181 3736 3185
rect 3776 3181 3780 3186
rect 4079 3180 4082 3280
rect 4173 3260 4177 3299
rect 4294 3298 4321 3299
rect 4339 3261 4343 3299
rect 4412 3276 4419 3299
rect 4079 3177 4165 3180
rect 4160 3161 4165 3177
rect 4174 3177 4178 3199
rect 4344 3188 4347 3201
rect 4270 3185 4347 3188
rect 4174 3173 4226 3177
rect 4048 3146 4096 3151
rect 3776 3120 3779 3127
rect 3776 3116 3800 3120
rect 3795 3080 3800 3116
rect 3908 3080 3912 3127
rect 3667 3075 3941 3080
rect 2981 3036 3424 3041
rect 4049 3026 4053 3146
rect 4180 3109 4185 3112
rect 4185 3066 4189 3108
rect 4223 3066 4226 3173
rect 4270 3066 4274 3185
rect 4413 3175 4419 3276
rect 4309 3172 4419 3175
rect 4487 3175 4492 3299
rect 4700 3211 4703 3311
rect 4794 3291 4798 3330
rect 4960 3292 4964 3330
rect 5033 3307 5040 3330
rect 4700 3208 4786 3211
rect 4558 3193 4565 3194
rect 4558 3186 4703 3193
rect 4781 3192 4786 3208
rect 4795 3208 4799 3230
rect 4965 3219 4968 3232
rect 4891 3216 4968 3219
rect 4795 3204 4847 3208
rect 4842 3203 4847 3204
rect 4309 3171 4347 3172
rect 4309 3167 4312 3171
rect 4352 3167 4356 3172
rect 4352 3106 4355 3113
rect 4352 3102 4376 3106
rect 4083 3061 4314 3066
rect 4371 3066 4376 3102
rect 4484 3066 4488 3113
rect 4322 3061 4517 3066
rect 4223 3060 4226 3061
rect 4558 3031 4565 3186
rect 4801 3140 4806 3143
rect 4806 3097 4810 3139
rect 4844 3098 4847 3203
rect 4704 3092 4843 3097
rect 4891 3097 4895 3216
rect 5034 3206 5040 3307
rect 4930 3203 5040 3206
rect 5108 3206 5113 3330
rect 4930 3202 4968 3203
rect 4930 3198 4933 3202
rect 4973 3198 4977 3203
rect 4973 3137 4976 3144
rect 4973 3133 4997 3137
rect 4992 3097 4997 3133
rect 5105 3120 5109 3144
rect 5105 3116 5110 3120
rect 5105 3097 5109 3116
rect 4853 3092 5138 3097
rect 1907 3021 2242 3025
rect 300 2948 332 2951
rect 1076 2949 1595 2955
rect 1076 2904 1082 2949
rect 75 2898 83 2902
rect 75 2797 79 2898
rect 371 2889 385 2893
rect 391 2889 392 2893
rect 163 2819 166 2886
rect 297 2869 353 2870
rect 297 2867 386 2869
rect 348 2866 386 2867
rect 468 2799 472 2896
rect 514 2889 528 2893
rect 534 2889 535 2893
rect 619 2821 624 2896
rect 677 2889 691 2893
rect 697 2889 698 2893
rect 618 2809 624 2821
rect 780 2828 785 2896
rect 833 2889 847 2893
rect 853 2889 854 2893
rect 937 2836 941 2895
rect 971 2889 985 2893
rect 991 2889 992 2893
rect 1114 2889 1128 2893
rect 1134 2889 1135 2893
rect 1216 2845 1221 2897
rect 1277 2889 1291 2893
rect 1297 2889 1298 2893
rect 1373 2856 1377 2896
rect 1433 2889 1447 2893
rect 1453 2889 1454 2893
rect 1859 2875 1863 2968
rect 1907 2962 1911 3021
rect 4049 3012 4054 3026
rect 2122 3008 4054 3012
rect 2122 2961 2126 3008
rect 4557 3003 4565 3031
rect 2433 3000 4565 3003
rect 2320 2995 4565 3000
rect 2320 2962 2325 2995
rect 2433 2994 4565 2995
rect 4557 2993 4565 2994
rect 1604 2871 1863 2875
rect 1604 2845 1609 2871
rect 1216 2841 1609 2845
rect 1604 2840 1609 2841
rect 937 2833 4669 2836
rect 937 2832 4614 2833
rect 4681 2833 4686 2836
rect 780 2824 784 2828
rect 780 2816 4066 2824
rect 618 2805 3458 2809
rect 620 2804 3458 2805
rect 75 2793 228 2797
rect 468 2796 2897 2799
rect 1389 2789 1838 2792
rect 301 2776 317 2781
rect 44 2754 282 2760
rect 312 2722 316 2776
rect 371 2740 385 2744
rect 391 2740 392 2744
rect 312 2720 355 2722
rect 312 2717 386 2720
rect 476 2671 481 2748
rect 514 2740 528 2744
rect 534 2740 535 2744
rect 614 2679 618 2748
rect 677 2740 691 2744
rect 697 2740 698 2744
rect 784 2688 788 2748
rect 833 2740 847 2744
rect 853 2740 854 2744
rect 938 2696 942 2748
rect 971 2740 985 2744
rect 991 2740 992 2744
rect 1082 2703 1085 2747
rect 1114 2740 1128 2744
rect 1134 2740 1135 2744
rect 1227 2710 1231 2748
rect 1389 2752 1392 2789
rect 1372 2748 1394 2752
rect 1527 2748 1816 2752
rect 1277 2740 1291 2744
rect 1297 2740 1298 2744
rect 1433 2740 1447 2744
rect 1453 2740 1454 2744
rect 1626 2710 1878 2712
rect 1227 2708 1878 2710
rect 1895 2710 1900 2711
rect 1227 2707 1635 2708
rect 1895 2706 1940 2710
rect 1895 2704 1900 2706
rect 1734 2703 1900 2704
rect 1082 2700 1900 2703
rect 1912 2696 1913 2697
rect 938 2693 1913 2696
rect 784 2684 1929 2688
rect 614 2676 1952 2679
rect 2383 2671 2387 2676
rect 2398 2671 2402 2676
rect 2413 2674 2417 2676
rect 2427 2674 2431 2676
rect 476 2668 1973 2671
rect 371 2615 385 2619
rect 391 2615 392 2619
rect 326 2595 339 2596
rect 326 2592 386 2595
rect 392 2592 395 2595
rect 469 2259 473 2623
rect 514 2615 528 2619
rect 534 2615 535 2619
rect 613 2313 618 2622
rect 677 2615 691 2619
rect 697 2615 698 2619
rect 779 2326 785 2622
rect 833 2615 847 2619
rect 853 2615 854 2619
rect 922 2335 927 2621
rect 971 2615 985 2619
rect 991 2615 992 2619
rect 1068 2461 1074 2622
rect 1114 2615 1128 2619
rect 1134 2615 1135 2619
rect 1222 2424 1227 2621
rect 1277 2615 1291 2619
rect 1297 2615 1298 2619
rect 1377 2398 1383 2620
rect 1433 2615 1447 2619
rect 1453 2615 1454 2619
rect 922 2331 1184 2335
rect 1969 2333 1973 2668
rect 2007 2411 2325 2414
rect 2007 2333 2012 2411
rect 2074 2367 2130 2371
rect 2135 2367 2136 2371
rect 779 2325 1011 2326
rect 781 2321 1011 2325
rect 613 2312 727 2313
rect 613 2306 863 2312
rect 705 2305 863 2306
rect 747 2259 767 2260
rect 469 2256 767 2259
rect 469 2255 753 2256
rect 858 2260 863 2305
rect 1004 2261 1010 2321
rect 773 2256 774 2260
rect 858 2256 910 2260
rect 858 2255 896 2256
rect 1004 2260 1054 2261
rect 916 2256 917 2260
rect 1004 2256 1073 2260
rect 1079 2256 1080 2260
rect 1180 2259 1183 2331
rect 1969 2330 2023 2333
rect 1969 2329 1983 2330
rect 1209 2259 1229 2260
rect 1180 2256 1229 2259
rect 1180 2255 1215 2256
rect 1235 2256 1236 2260
rect 1180 2254 1183 2255
rect 1980 1581 1983 2329
rect 2009 2257 2299 2260
rect 1997 2169 2004 2172
rect 2009 2172 2012 2257
rect 2076 2206 2132 2210
rect 2137 2206 2138 2210
rect 2009 2169 2025 2172
rect 1997 1648 2000 2169
rect 2007 2091 2042 2095
rect 2007 2018 2010 2091
rect 2075 2052 2131 2056
rect 2136 2052 2137 2056
rect 2007 2015 2015 2018
rect 2007 1715 2010 2015
rect 2020 2015 2024 2018
rect 2383 1943 2386 2671
rect 2398 2572 2401 2671
rect 2398 2538 2401 2567
rect 2413 2565 2416 2674
rect 2398 2159 2401 2533
rect 2015 1940 2386 1943
rect 2015 1872 2018 1940
rect 2075 1904 2131 1908
rect 2136 1904 2137 1908
rect 2020 1867 2024 1870
rect 2015 1781 2018 1865
rect 2015 1777 2077 1781
rect 2007 1711 2077 1715
rect 2270 1708 2294 1711
rect 1997 1644 2069 1648
rect 2270 1634 2274 1708
rect 2398 1648 2401 2154
rect 2413 2139 2416 2560
rect 2413 1692 2416 2134
rect 2427 2057 2430 2674
rect 2427 1797 2430 2052
rect 2537 1867 2566 1870
rect 2537 1812 2540 1867
rect 2427 1794 2568 1797
rect 2565 1786 2568 1794
rect 2565 1783 2612 1786
rect 2486 1692 2490 1701
rect 2413 1689 2469 1692
rect 2474 1689 2490 1692
rect 2496 1648 2500 1701
rect 2642 1648 2646 1782
rect 2398 1645 2646 1648
rect 2398 1631 2401 1645
rect 2350 1628 2401 1631
rect 1980 1577 2048 1581
<< m3contact >>
rect 365 3030 371 3035
rect 508 3030 514 3035
rect 671 3030 677 3035
rect 827 3030 833 3035
rect 965 3030 971 3035
rect 1108 3030 1114 3035
rect 1271 3030 1277 3035
rect 1427 3030 1433 3035
rect 365 2888 371 2893
rect 508 2888 514 2893
rect 671 2888 677 2893
rect 827 2888 833 2893
rect 965 2888 971 2893
rect 1108 2888 1114 2893
rect 1271 2888 1277 2893
rect 1427 2888 1433 2893
rect 365 2740 371 2746
rect 508 2739 514 2744
rect 671 2739 677 2744
rect 827 2739 833 2744
rect 965 2739 971 2744
rect 1108 2739 1114 2744
rect 1838 2787 1845 2792
rect 1816 2746 1823 2754
rect 1271 2739 1277 2744
rect 1427 2739 1433 2744
rect 1878 2708 1885 2715
rect 1940 2705 1948 2712
rect 1913 2693 1921 2700
rect 1929 2683 1936 2690
rect 1952 2675 1958 2680
rect 365 2614 371 2619
rect 508 2614 514 2619
rect 671 2614 677 2619
rect 827 2614 833 2619
rect 965 2614 971 2619
rect 1108 2614 1114 2619
rect 1271 2614 1277 2619
rect 1427 2614 1433 2619
rect 2325 2409 2330 2414
rect 2004 2169 2009 2174
rect 2015 2013 2020 2019
rect 2014 1865 2020 1872
<< m123contact >>
rect 2123 2697 2128 2702
rect 2131 2654 2136 2659
rect 2122 2631 2127 2636
rect 2131 2588 2136 2593
rect 2122 2564 2127 2569
rect 2131 2521 2136 2526
rect 2122 2497 2127 2502
rect 2131 2454 2136 2459
rect 2122 2391 2127 2396
rect 1940 2298 1946 2304
rect 1876 2131 1884 2139
rect 1943 2133 1951 2141
rect 1838 1979 1845 1986
rect 1942 1979 1951 1986
rect 2131 2308 2136 2313
rect 2122 2230 2127 2235
rect 2157 2230 2162 2235
rect 2132 2188 2137 2193
rect 2007 2126 2014 2133
rect 2122 2076 2127 2081
rect 2131 2034 2136 2039
rect 2017 1972 2023 1978
rect 2122 1928 2127 1933
rect 2131 1886 2136 1891
rect 2028 1818 2034 1824
rect 2122 1802 2127 1807
rect 2131 1759 2136 1764
rect 2122 1736 2127 1741
rect 2131 1693 2136 1698
rect 2122 1669 2127 1674
rect 2383 1706 2388 1711
rect 2384 1673 2389 1678
rect 2783 2507 2788 2512
rect 2730 2180 2735 2185
rect 2808 2118 2813 2123
rect 2834 1854 2839 1859
rect 2435 1781 2440 1786
rect 2131 1626 2136 1631
rect 2122 1602 2127 1607
rect 2131 1559 2136 1564
<< metal3 >>
rect 366 2893 370 3030
rect 509 2893 513 3030
rect 672 2893 676 3030
rect 828 2893 832 3030
rect 966 2893 970 3030
rect 1109 2893 1113 3030
rect 1272 2893 1276 3030
rect 1428 2893 1432 3030
rect 366 2746 370 2888
rect 509 2744 513 2888
rect 672 2744 676 2888
rect 828 2744 832 2888
rect 966 2744 970 2888
rect 1109 2744 1113 2888
rect 1272 2744 1276 2888
rect 1428 2744 1432 2888
rect 366 2619 370 2740
rect 509 2619 513 2739
rect 672 2619 676 2739
rect 828 2619 832 2739
rect 966 2726 970 2739
rect 965 2722 970 2726
rect 965 2670 969 2722
rect 965 2666 970 2670
rect 966 2619 970 2666
rect 1109 2619 1113 2739
rect 1272 2725 1276 2739
rect 1271 2714 1276 2725
rect 1428 2722 1432 2739
rect 1427 2714 1432 2722
rect 1271 2670 1275 2714
rect 1427 2670 1431 2714
rect 1271 2665 1276 2670
rect 1272 2619 1276 2665
rect 1427 2662 1432 2670
rect 1428 2619 1432 2662
rect 366 2587 370 2614
rect 509 2587 513 2614
rect 672 2587 676 2614
rect 828 2588 832 2614
rect 966 2597 970 2614
rect 1109 2589 1113 2614
rect 1272 2589 1276 2614
rect 1428 2589 1432 2614
rect 1817 1824 1821 2746
rect 1839 1986 1843 2787
rect 1879 2145 1883 2708
rect 1878 2139 1883 2145
rect 1913 1871 1918 2693
rect 1930 2018 1935 2683
rect 1940 2304 1944 2705
rect 1953 2172 1957 2675
rect 2123 2636 2127 2697
rect 2123 2569 2127 2631
rect 2123 2502 2127 2564
rect 2123 2396 2127 2497
rect 2123 2235 2127 2391
rect 1953 2169 2004 2172
rect 1951 2135 2012 2139
rect 2007 2133 2012 2135
rect 2123 2081 2127 2230
rect 1930 2015 2015 2018
rect 1941 1980 1942 1984
rect 1951 1980 2020 1984
rect 2017 1978 2020 1980
rect 2123 1933 2127 2076
rect 1913 1866 2014 1871
rect 2020 1866 2022 1871
rect 1817 1821 2028 1824
rect 2123 1807 2127 1928
rect 2123 1741 2127 1802
rect 2123 1674 2127 1736
rect 2123 1607 2127 1669
rect 2131 2593 2135 2654
rect 2131 2526 2135 2588
rect 2131 2459 2135 2521
rect 2131 2313 2135 2454
rect 2784 2414 2788 2507
rect 2330 2410 2788 2414
rect 2131 2193 2135 2308
rect 2162 2231 2730 2235
rect 2131 2188 2132 2193
rect 2131 2039 2135 2188
rect 2726 2182 2730 2231
rect 2131 2021 2135 2034
rect 2809 2021 2813 2118
rect 2131 2018 2813 2021
rect 2131 1891 2135 2018
rect 2131 1764 2135 1886
rect 2384 1783 2435 1786
rect 2131 1698 2135 1759
rect 2384 1711 2387 1783
rect 2131 1631 2135 1693
rect 2835 1678 2839 1854
rect 2389 1674 2839 1678
rect 2131 1564 2135 1626
<< labels >>
rlabel metal1 3381 3144 3381 3148 1 sub4
rlabel polysilicon 3163 3285 3166 3285 1 sub3
rlabel polysilicon 3726 3288 3729 3288 1 sub2
rlabel polysilicon 4302 3274 4305 3274 1 sub1
rlabel polysilicon 4923 3313 4926 3313 1 sub0
rlabel m2contact 2323 2958 2323 2959 1 gbu0
rlabel m2contact 2125 2957 2125 2958 1 gbu1
rlabel m2contact 1910 2958 1910 2959 1 gbu2
rlabel m2contact 1715 2957 1715 2958 1 gbu3
rlabel metal1 302 2799 302 2803 1 d1
rlabel metal1 1526 2897 1526 2901 7 goutb0
rlabel metal1 1064 3039 1064 3043 1 foutb3
rlabel polysilicon 406 3585 409 3585 1 sum3
rlabel polysilicon 969 3588 972 3588 1 sum2
rlabel polysilicon 1545 3574 1548 3574 1 sum1
rlabel polysilicon 2166 3613 2169 3613 1 sum0
rlabel metal1 624 3444 624 3448 1 sum4
rlabel metal1 1308 2264 1308 2268 1 and0
rlabel metal1 1152 2264 1152 2268 1 and1
rlabel metal1 989 2264 989 2268 1 and2
rlabel metal1 846 2264 846 2268 1 and3
rlabel metal1 916 2623 916 2627 1 iouta0
rlabel metal1 1207 2623 1207 2627 1 ioutb2
rlabel metal1 159 2888 159 2888 1 d3
rlabel metal1 1526 2623 1526 2627 7 ioutb0
rlabel metal1 1370 2623 1370 2627 1 ioutb1
rlabel metal1 1064 2623 1064 2627 1 ioutb3
rlabel metal1 770 2623 770 2627 1 iouta1
rlabel metal1 607 2623 607 2627 1 iouta2
rlabel metal1 464 2623 464 2627 1 iouta3
rlabel m2contact 1526 2748 1526 2752 7 houtb0
rlabel m2contact 1370 2748 1370 2752 1 houtb1
rlabel metal1 1207 2748 1207 2752 1 houtb2
rlabel metal1 1064 2748 1064 2752 1 houtb3
rlabel metal1 926 2748 926 2752 1 houta0
rlabel metal1 770 2748 770 2752 1 houta1
rlabel metal1 607 2748 607 2752 1 houta2
rlabel metal1 464 2748 464 2752 1 houta3
rlabel m2contact 298 2971 298 2975 1 d2
rlabel metal1 1370 2897 1370 2901 1 goutb1
rlabel metal1 1207 2897 1207 2901 1 goutb2
rlabel metal1 1064 2897 1064 2901 1 goutb3
rlabel metal1 926 2897 926 2901 1 gouta0
rlabel metal1 770 2897 770 2901 1 gouta1
rlabel metal1 607 2897 607 2901 1 gouta2
rlabel metal1 464 2897 464 2901 1 gouta3
rlabel metal1 1526 3039 1526 3043 7 foutb0
rlabel metal3 1430 3016 1430 3016 1 b0
rlabel metal1 1370 3039 1370 3043 1 foutb1
rlabel metal3 1274 3021 1274 3021 1 b1
rlabel metal3 1111 3019 1111 3019 1 b2
rlabel metal1 1207 3039 1207 3043 1 foutb2
rlabel metal3 968 3020 968 3020 1 b3
rlabel metal1 926 3039 926 3043 7 fouta0
rlabel metal3 830 3017 830 3017 1 a0
rlabel metal1 770 3039 770 3043 7 fouta1
rlabel metal3 674 3016 674 3016 1 a1
rlabel metal1 464 3039 464 3043 1 fouta3
rlabel metal1 607 3039 607 3043 7 fouta2
rlabel metal3 511 3019 511 3019 1 a2
rlabel metal1 425 3040 425 3040 1 outn
rlabel metal3 368 3010 368 3010 1 a3
rlabel metal1 143 2839 143 2839 1 S1
rlabel metal1 171 2922 171 2922 1 S0
rlabel metal1 296 2890 296 2894 1 d0
rlabel metal1 192 2905 192 2905 1 gnd
rlabel metal1 185 2944 185 2944 4 vdd
rlabel metal3 368 2758 368 2758 1 chi
rlabel metal1 2883 1897 2883 1901 1 l
rlabel metal1 2892 2677 2892 2681 1 g
rlabel metal1 2961 2149 2961 2153 1 e
<< end >>
