magic
tech scmos
timestamp 1700138227
<< nwell >>
rect -410 -258 -374 -239
rect -367 -258 -340 -239
rect -458 -309 -433 -292
rect -546 -342 -511 -323
rect -504 -342 -477 -323
rect -413 -339 -375 -320
rect -368 -339 -341 -320
rect -458 -392 -433 -375
rect -409 -428 -373 -409
rect -366 -410 -341 -409
rect -366 -428 -339 -410
<< ntransistor >>
rect -398 -282 -396 -277
rect -389 -282 -387 -277
rect -356 -282 -354 -277
rect -446 -326 -444 -322
rect -535 -366 -533 -361
rect -526 -366 -524 -361
rect -493 -366 -491 -361
rect -399 -363 -397 -358
rect -390 -363 -388 -358
rect -357 -363 -355 -358
rect -446 -408 -444 -404
rect -397 -452 -395 -447
rect -388 -452 -386 -447
rect -355 -452 -353 -447
<< ptransistor >>
rect -398 -251 -396 -246
rect -389 -251 -387 -246
rect -356 -251 -354 -246
rect -446 -303 -444 -299
rect -535 -335 -533 -330
rect -526 -335 -524 -330
rect -493 -335 -491 -330
rect -399 -332 -397 -327
rect -390 -332 -388 -327
rect -357 -332 -355 -327
rect -446 -386 -444 -382
rect -397 -421 -395 -416
rect -388 -421 -386 -416
rect -355 -421 -353 -416
<< ndiffusion >>
rect -403 -278 -398 -277
rect -399 -282 -398 -278
rect -396 -282 -389 -277
rect -387 -281 -385 -277
rect -387 -282 -381 -281
rect -361 -279 -356 -277
rect -357 -282 -356 -279
rect -354 -280 -351 -277
rect -354 -282 -347 -280
rect -447 -326 -446 -322
rect -444 -326 -443 -322
rect -540 -362 -535 -361
rect -536 -366 -535 -362
rect -533 -366 -526 -361
rect -524 -365 -522 -361
rect -524 -366 -518 -365
rect -498 -363 -493 -361
rect -494 -366 -493 -363
rect -491 -364 -488 -361
rect -491 -366 -484 -364
rect -404 -359 -399 -358
rect -400 -363 -399 -359
rect -397 -363 -390 -358
rect -388 -362 -386 -358
rect -388 -363 -382 -362
rect -362 -360 -357 -358
rect -358 -363 -357 -360
rect -355 -361 -352 -358
rect -355 -363 -348 -361
rect -447 -408 -446 -404
rect -444 -408 -443 -404
rect -402 -448 -397 -447
rect -398 -452 -397 -448
rect -395 -452 -388 -447
rect -386 -451 -384 -447
rect -386 -452 -380 -451
rect -360 -449 -355 -447
rect -356 -452 -355 -449
rect -353 -450 -350 -447
rect -353 -452 -346 -450
<< pdiffusion >>
rect -399 -249 -398 -246
rect -403 -251 -398 -249
rect -396 -248 -389 -246
rect -396 -251 -394 -248
rect -390 -251 -389 -248
rect -387 -249 -385 -246
rect -387 -251 -381 -249
rect -357 -249 -356 -246
rect -361 -251 -356 -249
rect -354 -250 -351 -246
rect -354 -251 -347 -250
rect -447 -303 -446 -299
rect -444 -303 -443 -299
rect -536 -333 -535 -330
rect -540 -335 -535 -333
rect -533 -332 -526 -330
rect -533 -335 -531 -332
rect -527 -335 -526 -332
rect -524 -333 -522 -330
rect -524 -335 -518 -333
rect -494 -333 -493 -330
rect -498 -335 -493 -333
rect -491 -334 -488 -330
rect -491 -335 -484 -334
rect -400 -330 -399 -327
rect -404 -332 -399 -330
rect -397 -329 -390 -327
rect -397 -332 -395 -329
rect -391 -332 -390 -329
rect -388 -330 -386 -327
rect -388 -332 -382 -330
rect -358 -330 -357 -327
rect -362 -332 -357 -330
rect -355 -331 -352 -327
rect -355 -332 -348 -331
rect -447 -386 -446 -382
rect -444 -386 -443 -382
rect -398 -419 -397 -416
rect -402 -421 -397 -419
rect -395 -418 -388 -416
rect -395 -421 -393 -418
rect -389 -421 -388 -418
rect -386 -419 -384 -416
rect -386 -421 -380 -419
rect -356 -419 -355 -416
rect -360 -421 -355 -419
rect -353 -420 -350 -416
rect -353 -421 -346 -420
<< ndcontact >>
rect -403 -282 -399 -278
rect -385 -281 -381 -277
rect -361 -283 -357 -279
rect -351 -280 -347 -276
rect -451 -326 -447 -322
rect -443 -326 -439 -322
rect -540 -366 -536 -362
rect -522 -365 -518 -361
rect -498 -367 -494 -363
rect -488 -364 -484 -360
rect -404 -363 -400 -359
rect -386 -362 -382 -358
rect -362 -364 -358 -360
rect -352 -361 -348 -357
rect -451 -408 -447 -404
rect -443 -408 -439 -404
rect -402 -452 -398 -448
rect -384 -451 -380 -447
rect -360 -453 -356 -449
rect -350 -450 -346 -446
<< pdcontact >>
rect -403 -249 -399 -245
rect -394 -252 -390 -248
rect -385 -249 -381 -245
rect -361 -249 -357 -245
rect -351 -250 -347 -246
rect -451 -303 -447 -299
rect -443 -303 -439 -299
rect -540 -333 -536 -329
rect -531 -336 -527 -332
rect -522 -333 -518 -329
rect -498 -333 -494 -329
rect -488 -334 -484 -330
rect -404 -330 -400 -326
rect -395 -333 -391 -329
rect -386 -330 -382 -326
rect -362 -330 -358 -326
rect -352 -331 -348 -327
rect -451 -386 -447 -382
rect -443 -386 -439 -382
rect -402 -419 -398 -415
rect -393 -422 -389 -418
rect -384 -419 -380 -415
rect -360 -419 -356 -415
rect -350 -420 -346 -416
<< polysilicon >>
rect -461 -242 -410 -239
rect -582 -288 -471 -285
rect -582 -373 -578 -288
rect -461 -292 -457 -242
rect -339 -242 -331 -239
rect -398 -246 -396 -243
rect -389 -246 -387 -243
rect -398 -261 -396 -251
rect -356 -246 -354 -243
rect -397 -265 -396 -261
rect -398 -277 -396 -265
rect -389 -270 -387 -251
rect -356 -262 -354 -251
rect -355 -266 -354 -262
rect -388 -274 -387 -270
rect -389 -277 -387 -274
rect -356 -277 -354 -266
rect -398 -285 -396 -282
rect -389 -285 -387 -282
rect -356 -285 -354 -282
rect -446 -288 -412 -286
rect -461 -295 -460 -292
rect -431 -296 -409 -293
rect -446 -299 -444 -296
rect -446 -313 -444 -303
rect -450 -315 -444 -313
rect -446 -322 -444 -315
rect -413 -320 -409 -296
rect -335 -320 -331 -242
rect -476 -326 -467 -323
rect -339 -324 -331 -320
rect -535 -330 -533 -327
rect -526 -330 -524 -327
rect -535 -345 -533 -335
rect -493 -330 -491 -327
rect -534 -349 -533 -345
rect -535 -361 -533 -349
rect -526 -354 -524 -335
rect -493 -346 -491 -335
rect -492 -350 -491 -346
rect -525 -358 -524 -354
rect -526 -361 -524 -358
rect -493 -361 -491 -350
rect -535 -369 -533 -366
rect -526 -369 -524 -366
rect -493 -369 -491 -366
rect -582 -376 -547 -373
rect -482 -412 -479 -377
rect -470 -375 -467 -326
rect -446 -329 -444 -326
rect -399 -327 -397 -324
rect -390 -327 -388 -324
rect -434 -360 -431 -334
rect -399 -342 -397 -332
rect -357 -327 -355 -324
rect -398 -346 -397 -342
rect -399 -358 -397 -346
rect -390 -351 -388 -332
rect -357 -343 -355 -332
rect -356 -347 -355 -343
rect -389 -355 -388 -351
rect -390 -358 -388 -355
rect -357 -358 -355 -347
rect -434 -363 -407 -360
rect -410 -367 -407 -363
rect -399 -366 -397 -363
rect -390 -366 -388 -363
rect -357 -366 -355 -363
rect -470 -378 -460 -375
rect -430 -378 -405 -375
rect -446 -382 -444 -379
rect -466 -412 -463 -392
rect -446 -396 -444 -386
rect -450 -398 -444 -396
rect -446 -404 -444 -398
rect -446 -411 -444 -408
rect -409 -409 -405 -378
rect -335 -409 -331 -324
rect -482 -415 -459 -412
rect -337 -412 -331 -409
rect -435 -456 -432 -416
rect -397 -416 -395 -413
rect -388 -416 -386 -413
rect -397 -431 -395 -421
rect -355 -416 -353 -413
rect -396 -435 -395 -431
rect -397 -447 -395 -435
rect -388 -440 -386 -421
rect -355 -432 -353 -421
rect -354 -436 -353 -432
rect -387 -444 -386 -440
rect -388 -447 -386 -444
rect -355 -447 -353 -436
rect -397 -455 -395 -452
rect -388 -455 -386 -452
rect -355 -455 -353 -452
rect -435 -459 -409 -456
<< polycontact >>
rect -471 -289 -467 -285
rect -410 -243 -406 -239
rect -343 -243 -339 -239
rect -401 -265 -397 -261
rect -359 -266 -355 -262
rect -392 -274 -388 -270
rect -450 -289 -446 -285
rect -412 -289 -408 -285
rect -460 -296 -456 -292
rect -435 -296 -431 -292
rect -454 -316 -450 -312
rect -480 -327 -476 -323
rect -413 -324 -409 -320
rect -343 -324 -339 -320
rect -538 -349 -534 -345
rect -496 -350 -492 -346
rect -529 -358 -525 -354
rect -547 -377 -543 -373
rect -483 -377 -479 -373
rect -435 -334 -431 -330
rect -402 -346 -398 -342
rect -360 -347 -356 -343
rect -393 -355 -389 -351
rect -410 -371 -406 -367
rect -460 -379 -456 -375
rect -434 -379 -430 -375
rect -467 -392 -463 -388
rect -454 -399 -450 -395
rect -459 -416 -455 -412
rect -436 -416 -432 -412
rect -409 -413 -405 -409
rect -341 -413 -337 -409
rect -400 -435 -396 -431
rect -358 -436 -354 -432
rect -391 -444 -387 -440
rect -409 -460 -405 -456
<< metal1 >>
rect -406 -242 -343 -239
rect -403 -245 -399 -242
rect -385 -245 -381 -242
rect -361 -245 -357 -242
rect -572 -265 -401 -261
rect -394 -262 -390 -252
rect -351 -262 -347 -250
rect -572 -363 -568 -265
rect -394 -266 -359 -262
rect -351 -266 -343 -262
rect -424 -274 -392 -270
rect -467 -288 -450 -285
rect -456 -295 -435 -292
rect -450 -299 -447 -295
rect -443 -312 -439 -303
rect -424 -312 -420 -274
rect -385 -277 -381 -266
rect -351 -276 -347 -266
rect -403 -286 -399 -282
rect -361 -286 -357 -283
rect -408 -289 -343 -286
rect -555 -316 -454 -312
rect -443 -316 -420 -312
rect -555 -335 -551 -316
rect -443 -322 -439 -316
rect -545 -326 -480 -323
rect -540 -329 -536 -326
rect -522 -329 -518 -326
rect -552 -340 -551 -335
rect -555 -345 -551 -340
rect -498 -329 -494 -326
rect -450 -330 -447 -326
rect -555 -349 -538 -345
rect -531 -346 -527 -336
rect -488 -346 -484 -334
rect -466 -333 -435 -330
rect -531 -350 -496 -346
rect -488 -350 -480 -346
rect -555 -358 -529 -354
rect -555 -363 -551 -358
rect -522 -361 -518 -350
rect -572 -367 -551 -363
rect -555 -395 -551 -367
rect -488 -360 -484 -350
rect -540 -373 -536 -366
rect -498 -373 -494 -367
rect -543 -376 -483 -373
rect -466 -388 -463 -333
rect -424 -342 -420 -316
rect -409 -323 -343 -320
rect -404 -326 -400 -323
rect -386 -326 -382 -323
rect -362 -326 -358 -323
rect -424 -346 -402 -342
rect -395 -343 -391 -333
rect -352 -343 -348 -331
rect -395 -347 -360 -343
rect -352 -347 -344 -343
rect -418 -355 -393 -351
rect -456 -378 -434 -375
rect -450 -382 -447 -378
rect -443 -395 -439 -386
rect -418 -395 -414 -355
rect -386 -358 -382 -347
rect -352 -357 -348 -347
rect -404 -367 -400 -363
rect -362 -367 -358 -364
rect -406 -370 -344 -367
rect -555 -399 -454 -395
rect -443 -399 -414 -395
rect -443 -404 -439 -399
rect -450 -412 -447 -408
rect -455 -415 -436 -412
rect -425 -431 -421 -399
rect -405 -412 -341 -409
rect -402 -415 -398 -412
rect -384 -415 -380 -412
rect -360 -415 -356 -412
rect -425 -435 -400 -431
rect -393 -432 -389 -422
rect -350 -432 -346 -420
rect -393 -436 -358 -432
rect -350 -436 -342 -432
rect -406 -444 -391 -440
rect -384 -447 -380 -436
rect -350 -446 -346 -436
rect -402 -456 -398 -452
rect -360 -456 -356 -453
rect -405 -459 -342 -456
<< m2contact >>
rect -557 -340 -552 -335
rect -411 -445 -406 -440
<< metal2 >>
rect -565 -339 -557 -335
rect -565 -440 -561 -339
rect -565 -444 -411 -440
<< labels >>
rlabel metal1 -455 -293 -455 -293 4 vdd
rlabel metal1 -448 -332 -448 -332 1 gnd
rlabel metal1 -344 -347 -344 -343 1 d0
rlabel metal1 -343 -266 -343 -262 1 d2
rlabel metal1 -480 -350 -480 -346 1 d3
rlabel metal1 -342 -436 -342 -432 1 d1
rlabel metal1 -469 -315 -469 -315 1 S0
rlabel metal1 -497 -398 -497 -398 1 S1
<< end >>
