magic
tech scmos
timestamp 1698905099
<< nwell >>
rect -13 7 12 24
<< ntransistor >>
rect -1 -10 1 -6
<< ptransistor >>
rect -1 13 1 17
<< ndiffusion >>
rect -2 -10 -1 -6
rect 1 -10 2 -6
<< pdiffusion >>
rect -2 13 -1 17
rect 1 13 2 17
<< ndcontact >>
rect -6 -10 -2 -6
rect 2 -10 6 -6
<< pdcontact >>
rect -6 13 -2 17
rect 2 13 6 17
<< polysilicon >>
rect -1 17 1 20
rect -1 3 1 13
rect -5 1 1 3
rect -1 -6 1 1
rect -1 -13 1 -10
<< polycontact >>
rect -9 0 -5 4
<< metal1 >>
rect -13 21 12 24
rect -5 17 -2 21
rect 2 4 6 13
rect -12 0 -9 4
rect 2 0 9 4
rect 2 -6 6 0
rect -5 -14 -2 -10
rect -12 -17 12 -14
<< labels >>
rlabel metal1 -12 0 -12 4 3 in
rlabel metal1 9 0 9 4 7 out
rlabel metal1 -3 -16 -3 -16 1 gnd
rlabel metal1 -10 23 -10 23 4 vdd
<< end >>
