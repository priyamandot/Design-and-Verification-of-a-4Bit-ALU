magic
tech scmos
timestamp 1700302574
<< nwell >>
rect 0 90 55 109
rect 63 90 90 109
<< ntransistor >>
rect 11 66 13 71
rect 20 66 22 71
rect 29 66 31 71
rect 38 66 40 71
rect 74 66 76 71
<< ptransistor >>
rect 11 97 13 102
rect 20 97 22 102
rect 29 97 31 102
rect 38 97 40 102
rect 74 97 76 102
<< ndiffusion >>
rect 6 70 11 71
rect 10 66 11 70
rect 13 66 20 71
rect 22 66 29 71
rect 31 66 38 71
rect 40 66 42 71
rect 46 66 51 71
rect 69 69 74 71
rect 73 66 74 69
rect 76 68 79 71
rect 76 66 83 68
<< pdiffusion >>
rect 10 99 11 102
rect 6 97 11 99
rect 13 100 20 102
rect 13 97 15 100
rect 19 97 20 100
rect 22 99 24 102
rect 28 99 29 102
rect 22 97 29 99
rect 31 100 38 102
rect 31 97 33 100
rect 37 97 38 100
rect 40 99 42 102
rect 40 97 46 99
rect 73 99 74 102
rect 69 97 74 99
rect 76 98 79 102
rect 76 97 83 98
<< ndcontact >>
rect 6 66 10 70
rect 42 66 46 72
rect 69 65 73 69
rect 79 68 83 72
<< pdcontact >>
rect 6 99 10 103
rect 15 96 19 100
rect 24 99 28 103
rect 33 96 37 100
rect 42 99 46 103
rect 69 99 73 103
rect 79 98 83 102
<< polysilicon >>
rect 11 102 13 105
rect 20 102 22 105
rect 11 71 13 97
rect 29 102 31 105
rect 38 102 40 105
rect 20 71 22 97
rect 29 71 31 97
rect 74 102 76 105
rect 38 71 40 97
rect 74 86 76 97
rect 75 82 76 86
rect 74 71 76 82
rect 11 63 13 66
rect 20 63 22 66
rect 29 63 31 66
rect 38 63 40 66
rect 74 63 76 66
<< polycontact >>
rect 71 82 75 86
<< metal1 >>
rect 1 106 87 109
rect 6 103 10 106
rect 24 103 28 106
rect 42 103 46 106
rect 15 86 19 96
rect 69 103 73 106
rect 33 86 37 96
rect 79 86 83 98
rect 15 82 71 86
rect 79 82 87 86
rect 42 72 46 82
rect 79 72 83 82
rect 6 62 10 66
rect 69 62 73 65
rect 1 59 87 62
<< labels >>
rlabel metal1 24 60 24 60 1 gnd
rlabel metal1 38 108 38 108 5 vdd
rlabel polysilicon 12 83 12 83 1 A
rlabel polysilicon 21 80 21 80 1 B
rlabel polysilicon 30 80 30 80 1 C
rlabel polysilicon 39 80 39 80 1 D
rlabel metal1 87 82 87 86 7 out
<< end >>
