magic
tech scmos
timestamp 1700141014
<< nwell >>
rect 575 80 610 99
rect 617 80 644 99
rect 680 80 715 99
rect 722 80 749 99
rect 785 80 820 99
rect 827 80 854 99
rect 879 80 914 99
rect 921 80 948 99
rect 974 80 1009 99
rect 1016 80 1043 99
rect 1072 80 1107 99
rect 1114 80 1141 99
rect 1170 80 1205 99
rect 1212 80 1239 99
rect 1265 80 1300 99
rect 1307 80 1334 99
<< ntransistor >>
rect 586 56 588 61
rect 595 56 597 61
rect 628 56 630 61
rect 691 56 693 61
rect 700 56 702 61
rect 733 56 735 61
rect 796 56 798 61
rect 805 56 807 61
rect 838 56 840 61
rect 890 56 892 61
rect 899 56 901 61
rect 932 56 934 61
rect 985 56 987 61
rect 994 56 996 61
rect 1027 56 1029 61
rect 1083 56 1085 61
rect 1092 56 1094 61
rect 1125 56 1127 61
rect 1181 56 1183 61
rect 1190 56 1192 61
rect 1223 56 1225 61
rect 1276 56 1278 61
rect 1285 56 1287 61
rect 1318 56 1320 61
<< ptransistor >>
rect 586 87 588 92
rect 595 87 597 92
rect 628 87 630 92
rect 691 87 693 92
rect 700 87 702 92
rect 733 87 735 92
rect 796 87 798 92
rect 805 87 807 92
rect 838 87 840 92
rect 890 87 892 92
rect 899 87 901 92
rect 932 87 934 92
rect 985 87 987 92
rect 994 87 996 92
rect 1027 87 1029 92
rect 1083 87 1085 92
rect 1092 87 1094 92
rect 1125 87 1127 92
rect 1181 87 1183 92
rect 1190 87 1192 92
rect 1223 87 1225 92
rect 1276 87 1278 92
rect 1285 87 1287 92
rect 1318 87 1320 92
<< ndiffusion >>
rect 581 60 586 61
rect 585 56 586 60
rect 588 56 595 61
rect 597 57 598 61
rect 597 56 602 57
rect 623 59 628 61
rect 627 56 628 59
rect 630 58 633 61
rect 630 56 637 58
rect 686 60 691 61
rect 690 56 691 60
rect 693 56 700 61
rect 702 57 703 61
rect 702 56 707 57
rect 728 59 733 61
rect 732 56 733 59
rect 735 58 738 61
rect 735 56 742 58
rect 791 60 796 61
rect 795 56 796 60
rect 798 56 805 61
rect 807 57 808 61
rect 807 56 812 57
rect 833 59 838 61
rect 837 56 838 59
rect 840 58 843 61
rect 840 56 847 58
rect 885 60 890 61
rect 889 56 890 60
rect 892 56 899 61
rect 901 57 902 61
rect 901 56 906 57
rect 927 59 932 61
rect 931 56 932 59
rect 934 58 937 61
rect 934 56 941 58
rect 980 60 985 61
rect 984 56 985 60
rect 987 56 994 61
rect 996 57 997 61
rect 996 56 1001 57
rect 1022 59 1027 61
rect 1026 56 1027 59
rect 1029 58 1032 61
rect 1029 56 1036 58
rect 1078 60 1083 61
rect 1082 56 1083 60
rect 1085 56 1092 61
rect 1094 57 1095 61
rect 1094 56 1099 57
rect 1120 59 1125 61
rect 1124 56 1125 59
rect 1127 58 1130 61
rect 1127 56 1134 58
rect 1176 60 1181 61
rect 1180 56 1181 60
rect 1183 56 1190 61
rect 1192 57 1193 61
rect 1192 56 1197 57
rect 1218 59 1223 61
rect 1222 56 1223 59
rect 1225 58 1228 61
rect 1225 56 1232 58
rect 1271 60 1276 61
rect 1275 56 1276 60
rect 1278 56 1285 61
rect 1287 57 1288 61
rect 1287 56 1292 57
rect 1313 59 1318 61
rect 1317 56 1318 59
rect 1320 58 1323 61
rect 1320 56 1327 58
<< pdiffusion >>
rect 585 89 586 92
rect 581 87 586 89
rect 588 90 595 92
rect 588 87 590 90
rect 594 87 595 90
rect 597 89 599 92
rect 597 87 603 89
rect 627 89 628 92
rect 623 87 628 89
rect 630 88 633 92
rect 630 87 637 88
rect 690 89 691 92
rect 686 87 691 89
rect 693 90 700 92
rect 693 87 695 90
rect 699 87 700 90
rect 702 89 704 92
rect 702 87 708 89
rect 732 89 733 92
rect 728 87 733 89
rect 735 88 738 92
rect 735 87 742 88
rect 795 89 796 92
rect 791 87 796 89
rect 798 90 805 92
rect 798 87 800 90
rect 804 87 805 90
rect 807 89 809 92
rect 807 87 813 89
rect 837 89 838 92
rect 833 87 838 89
rect 840 88 843 92
rect 840 87 847 88
rect 889 89 890 92
rect 885 87 890 89
rect 892 90 899 92
rect 892 87 894 90
rect 898 87 899 90
rect 901 89 903 92
rect 901 87 907 89
rect 931 89 932 92
rect 927 87 932 89
rect 934 88 937 92
rect 934 87 941 88
rect 984 89 985 92
rect 980 87 985 89
rect 987 90 994 92
rect 987 87 989 90
rect 993 87 994 90
rect 996 89 998 92
rect 996 87 1002 89
rect 1026 89 1027 92
rect 1022 87 1027 89
rect 1029 88 1032 92
rect 1029 87 1036 88
rect 1082 89 1083 92
rect 1078 87 1083 89
rect 1085 90 1092 92
rect 1085 87 1087 90
rect 1091 87 1092 90
rect 1094 89 1096 92
rect 1094 87 1100 89
rect 1124 89 1125 92
rect 1120 87 1125 89
rect 1127 88 1130 92
rect 1127 87 1134 88
rect 1180 89 1181 92
rect 1176 87 1181 89
rect 1183 90 1190 92
rect 1183 87 1185 90
rect 1189 87 1190 90
rect 1192 89 1194 92
rect 1192 87 1198 89
rect 1222 89 1223 92
rect 1218 87 1223 89
rect 1225 88 1228 92
rect 1225 87 1232 88
rect 1275 89 1276 92
rect 1271 87 1276 89
rect 1278 90 1285 92
rect 1278 87 1280 90
rect 1284 87 1285 90
rect 1287 89 1289 92
rect 1287 87 1293 89
rect 1317 89 1318 92
rect 1313 87 1318 89
rect 1320 88 1323 92
rect 1320 87 1327 88
<< ndcontact >>
rect 581 56 585 60
rect 598 57 602 61
rect 623 55 627 59
rect 633 58 637 62
rect 686 56 690 60
rect 703 57 707 61
rect 728 55 732 59
rect 738 58 742 62
rect 791 56 795 60
rect 808 57 812 61
rect 833 55 837 59
rect 843 58 847 62
rect 885 56 889 60
rect 902 57 906 61
rect 927 55 931 59
rect 937 58 941 62
rect 980 56 984 60
rect 997 57 1001 61
rect 1022 55 1026 59
rect 1032 58 1036 62
rect 1078 56 1082 60
rect 1095 57 1099 61
rect 1120 55 1124 59
rect 1130 58 1134 62
rect 1176 56 1180 60
rect 1193 57 1197 61
rect 1218 55 1222 59
rect 1228 58 1232 62
rect 1271 56 1275 60
rect 1288 57 1292 61
rect 1313 55 1317 59
rect 1323 58 1327 62
<< pdcontact >>
rect 581 89 585 93
rect 590 86 594 90
rect 599 89 603 93
rect 623 89 627 93
rect 633 88 637 92
rect 686 89 690 93
rect 695 86 699 90
rect 704 89 708 93
rect 728 89 732 93
rect 738 88 742 92
rect 791 89 795 93
rect 800 86 804 90
rect 809 89 813 93
rect 833 89 837 93
rect 843 88 847 92
rect 885 89 889 93
rect 894 86 898 90
rect 903 89 907 93
rect 927 89 931 93
rect 937 88 941 92
rect 980 89 984 93
rect 989 86 993 90
rect 998 89 1002 93
rect 1022 89 1026 93
rect 1032 88 1036 92
rect 1078 89 1082 93
rect 1087 86 1091 90
rect 1096 89 1100 93
rect 1120 89 1124 93
rect 1130 88 1134 92
rect 1176 89 1180 93
rect 1185 86 1189 90
rect 1194 89 1198 93
rect 1218 89 1222 93
rect 1228 88 1232 92
rect 1271 89 1275 93
rect 1280 86 1284 90
rect 1289 89 1293 93
rect 1313 89 1317 93
rect 1323 88 1327 92
<< polysilicon >>
rect 586 92 588 95
rect 595 92 597 95
rect 586 61 588 87
rect 628 92 630 95
rect 691 92 693 95
rect 700 92 702 95
rect 595 61 597 87
rect 628 76 630 87
rect 629 72 630 76
rect 628 61 630 72
rect 586 53 588 56
rect 595 53 597 56
rect 691 61 693 87
rect 733 92 735 95
rect 796 92 798 95
rect 805 92 807 95
rect 700 61 702 87
rect 733 76 735 87
rect 734 72 735 76
rect 733 61 735 72
rect 628 53 630 56
rect 691 53 693 56
rect 700 53 702 56
rect 796 61 798 87
rect 838 92 840 95
rect 890 92 892 95
rect 899 92 901 95
rect 805 61 807 87
rect 838 76 840 87
rect 839 72 840 76
rect 838 61 840 72
rect 733 53 735 56
rect 796 53 798 56
rect 805 53 807 56
rect 890 61 892 87
rect 932 92 934 95
rect 985 92 987 95
rect 994 92 996 95
rect 899 61 901 87
rect 932 76 934 87
rect 933 72 934 76
rect 932 61 934 72
rect 838 53 840 56
rect 890 53 892 56
rect 899 53 901 56
rect 985 61 987 87
rect 1027 92 1029 95
rect 1083 92 1085 95
rect 1092 92 1094 95
rect 994 61 996 87
rect 1027 76 1029 87
rect 1028 72 1029 76
rect 1027 61 1029 72
rect 932 53 934 56
rect 985 53 987 56
rect 994 53 996 56
rect 1083 61 1085 87
rect 1125 92 1127 95
rect 1181 92 1183 95
rect 1190 92 1192 95
rect 1092 61 1094 87
rect 1125 76 1127 87
rect 1126 72 1127 76
rect 1125 61 1127 72
rect 1027 53 1029 56
rect 1083 53 1085 56
rect 1092 53 1094 56
rect 1181 61 1183 87
rect 1223 92 1225 95
rect 1276 92 1278 95
rect 1285 92 1287 95
rect 1190 61 1192 87
rect 1223 76 1225 87
rect 1224 72 1225 76
rect 1223 61 1225 72
rect 1125 53 1127 56
rect 1181 53 1183 56
rect 1190 53 1192 56
rect 1276 61 1278 87
rect 1318 92 1320 95
rect 1285 61 1287 87
rect 1318 76 1320 87
rect 1319 72 1320 76
rect 1318 61 1320 72
rect 1223 53 1225 56
rect 1276 53 1278 56
rect 1285 53 1287 56
rect 1318 53 1320 56
<< polycontact >>
rect 625 72 629 76
rect 730 72 734 76
rect 835 72 839 76
rect 929 72 933 76
rect 1024 72 1028 76
rect 1122 72 1126 76
rect 1220 72 1224 76
rect 1315 72 1319 76
<< metal1 >>
rect 576 96 1334 99
rect 581 93 585 96
rect 599 93 603 96
rect 623 93 627 96
rect 686 93 690 96
rect 590 76 594 86
rect 704 93 708 96
rect 633 76 637 88
rect 728 93 732 96
rect 791 93 795 96
rect 695 76 699 86
rect 809 93 813 96
rect 738 76 742 88
rect 833 93 837 96
rect 885 93 889 96
rect 800 76 804 86
rect 903 93 907 96
rect 843 76 847 88
rect 927 93 931 96
rect 980 93 984 96
rect 894 76 898 86
rect 998 93 1002 96
rect 937 76 941 88
rect 1022 93 1026 96
rect 1078 93 1082 96
rect 989 76 993 86
rect 1096 93 1100 96
rect 1032 76 1036 88
rect 1120 93 1124 96
rect 1176 93 1180 96
rect 1087 76 1091 86
rect 1194 93 1198 96
rect 1130 76 1134 88
rect 1218 93 1222 96
rect 1271 93 1275 96
rect 1185 76 1189 86
rect 1289 93 1293 96
rect 1228 76 1232 88
rect 1313 93 1317 96
rect 1280 76 1284 86
rect 1323 76 1327 88
rect 590 72 625 76
rect 633 72 641 76
rect 695 72 730 76
rect 738 72 746 76
rect 800 72 835 76
rect 843 72 851 76
rect 894 72 929 76
rect 937 72 945 76
rect 989 72 1024 76
rect 1032 72 1040 76
rect 1087 72 1122 76
rect 1130 72 1138 76
rect 1185 72 1220 76
rect 1228 72 1236 76
rect 1280 72 1315 76
rect 1323 72 1331 76
rect 598 61 602 72
rect 633 62 637 72
rect 581 52 585 56
rect 703 61 707 72
rect 623 52 627 55
rect 738 62 742 72
rect 686 52 690 56
rect 808 61 812 72
rect 728 52 732 55
rect 843 62 847 72
rect 791 52 795 56
rect 902 61 906 72
rect 833 52 837 55
rect 937 62 941 72
rect 885 52 889 56
rect 997 61 1001 72
rect 927 52 931 55
rect 1032 62 1036 72
rect 980 52 984 56
rect 1095 61 1099 72
rect 1022 52 1026 55
rect 1130 62 1134 72
rect 1078 52 1082 56
rect 1193 61 1197 72
rect 1120 52 1124 55
rect 1228 62 1232 72
rect 1176 52 1180 56
rect 1288 61 1292 72
rect 1218 52 1222 55
rect 1323 62 1327 72
rect 1271 52 1275 56
rect 1313 52 1317 55
rect 576 49 1331 52
<< end >>
